@Filename: c:\vsm-lv\Will\data\AJA335e-FePtFeRh_1030nm_Tann_6\AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_50deg.VHD
@Measurement Controlfilename: C:\vsm-lv\Will\Recipes\10kOe OoP loop 50deg.VHC
@Signal Manipulation filename: c:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA335e-FePtFeRh_1030nm_Tann_600C
@Date: 05 November 2019    (2019-05-11)
@Time: 13:12:43
@Test ID: AJA335e_FePt_FeRh_Pt_600deg_annealed_OoP_RT
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 90.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Sample Temperature to 50.0948 [degC] and wait 60.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Applied Field to 9999.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 3:      Set Auto Range Signal to 12.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 5
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 5.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 10000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To: 50.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: 50.0000 [Oe] To: -50.0000 [Oe] Min Stepsize/Sweeprate =  2.0000 [Oe] Max Stepsize/Sweeprate =  2.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -50.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -10000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 4 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 20 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.706
@Y Coils Correction Factor: 0.964
@Sample Shape Correction Factor: 0.919
@Coil Angle Alpha: 42.300
@Coil Angle Beta: -47.320
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
15000.000000   1.000000
15249.000000   1.000524
15499.000000   1.000702
15750.000000   1.001233
16000.000000   1.001406
16250.000000   1.001585
16499.000000   1.001758
16749.000000   1.001937
16999.000000   1.002110
17249.000000   1.001937
17499.000000   1.002289
17749.000000   1.002289
17999.000000   1.002289
18249.000000   1.002462
18499.000000   1.002462
18748.000000   1.002462
18999.000000   1.002462
19249.000000   1.002462
19499.000000   1.002642
19749.000000   1.002642
19999.000000   1.002462
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = No
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 25 October 2019  12:02:56
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 5
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 13:12:43
@@Data
New Section: Section 0: 
2.965800E+1   5.005001E+1   5.005001E+1   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -1.432004E-1   2.379320E-1   -2.434958E-4   -4.963771E-5   4.963771E-5   -2.434958E-4   2.485037E-4   -1.684779E+2   -7.847787E+1   
5.500600E+1   5.007339E+1   5.007339E+1   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -1.229950E-1   2.152087E-1   -2.162044E-4   -4.972642E-5   4.972642E-5   -2.162044E-4   2.218492E-4   -1.670474E+2   -7.704739E+1   
8.046900E+1   5.006259E+1   5.006259E+1   8.998000E+3   8.998000E+3   9.000000E+1   8.998000E+3   8.998000E+3   -1.172666E-1   2.018458E-1   -2.039597E-4   -4.522702E-5   4.522702E-5   -2.039597E-4   2.089140E-4   -1.674973E+2   -7.749726E+1   
1.056150E+2   5.004449E+1   5.004449E+1   8.498000E+3   8.498000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -1.006590E-1   1.802847E-1   -1.796496E-4   -4.341449E-5   4.341449E-5   -1.796496E-4   1.848210E-4   -1.664143E+2   -7.641426E+1   
1.318130E+2   5.001980E+1   5.001980E+1   7.999000E+3   7.999000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -8.756420E-2   1.614147E-1   -1.592640E-4   -4.076318E-5   4.076318E-5   -1.592640E-4   1.643978E-4   -1.656435E+2   -7.564350E+1   
1.572170E+2   5.005270E+1   5.005270E+1   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -7.412695E-2   1.403727E-1   -1.372520E-4   -3.694512E-5   3.694512E-5   -1.372520E-4   1.421375E-4   -1.649344E+2   -7.493437E+1   
1.820090E+2   5.002599E+1   5.002599E+1   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -6.332970E-2   1.250429E-1   -1.205925E-4   -3.490892E-5   3.490892E-5   -1.205925E-4   1.255436E-4   -1.638554E+2   -7.385542E+1   
2.073530E+2   5.003741E+1   5.003741E+1   6.498000E+3   6.498000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -4.774151E-2   1.045016E-1   -9.757683E-5   -3.300911E-5   3.300911E-5   -9.757683E-5   1.030089E-4   -1.613099E+2   -7.130992E+1   
2.326840E+2   5.002499E+1   5.002499E+1   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -3.525527E-2   8.703589E-2   -7.848201E-5   -3.082572E-5   3.082572E-5   -7.848201E-5   8.431875E-5   -1.585564E+2   -6.855638E+1   
2.580990E+2   5.001351E+1   5.001351E+1   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -2.401586E-2   6.917195E-2   -5.989869E-5   -2.745979E-5   2.745979E-5   -5.989869E-5   6.589304E-5   -1.553715E+2   -6.537151E+1   
2.836430E+2   5.003439E+1   5.003439E+1   4.997000E+3   4.997000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -1.220827E-2   5.223301E-2   -4.156653E-5   -2.511885E-5   2.511885E-5   -4.156653E-5   4.856679E-5   -1.488552E+2   -5.885523E+1   
3.092350E+2   5.003130E+1   5.003130E+1   4.498000E+3   4.498000E+3   9.000000E+1   4.498000E+3   4.498000E+3   3.239757E-4   3.390198E-2   -2.187970E-5   -2.240378E-5   2.240378E-5   -2.187970E-5   3.131534E-5   -1.343220E+2   -4.432196E+1   
3.351110E+2   5.002441E+1   5.002441E+1   3.999000E+3   3.999000E+3   9.000000E+1   3.999000E+3   3.999000E+3   1.246506E-2   1.734829E-2   -3.592275E-6   -2.056137E-5   2.056137E-5   -3.592275E-6   2.087281E-5   -9.991012E+1   -9.910119E+0   
3.605140E+2   5.003799E+1   5.003799E+1   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   2.264387E-2   -3.485179E-4   1.422649E-5   -1.652026E-5   1.652026E-5   1.422649E-5   2.180165E-5   -4.926648E+1   4.073352E+1   
3.858180E+2   5.004781E+1   5.004781E+1   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   3.602039E-2   -1.835948E-2   3.422682E-5   -1.463889E-5   1.463889E-5   3.422682E-5   3.722597E-5   -2.315651E+1   6.684349E+1   
4.116350E+2   5.005029E+1   5.005029E+1   2.498000E+3   2.498000E+3   9.000000E+1   2.498000E+3   2.498000E+3   4.677906E-2   -3.619005E-2   5.249120E-5   -1.093922E-5   1.093922E-5   5.249120E-5   5.361896E-5   -1.177201E+1   7.822799E+1   
4.374210E+2   5.003799E+1   5.003799E+1   1.999000E+3   1.999000E+3   9.000000E+1   1.999000E+3   1.999000E+3   6.085664E-2   -5.462785E-2   7.320296E-5   -9.297318E-6   9.297318E-6   7.320296E-5   7.379101E-5   -7.238235E+0   8.276177E+1   
4.712690E+2   5.001260E+1   5.001260E+1   1.949000E+3   1.949000E+3   9.000000E+1   1.949000E+3   1.949000E+3   6.339842E-2   -5.625324E-2   7.583301E-5   -1.011466E-5   1.011466E-5   7.583301E-5   7.650459E-5   -7.597312E+0   8.240269E+1   
4.935040E+2   5.004171E+1   5.004171E+1   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   6.204425E-2   -5.738007E-2   7.572969E-5   -8.376387E-6   8.376387E-6   7.572969E-5   7.619153E-5   -6.311774E+0   8.368823E+1   
5.157870E+2   5.004769E+1   5.004769E+1   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   6.545303E-2   -5.953500E-2   7.924064E-5   -9.488791E-6   9.488791E-6   7.924064E-5   7.980674E-5   -6.828457E+0   8.317154E+1   
5.381120E+2   5.003460E+1   5.003460E+1   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   6.591444E-2   -6.091464E-2   8.042445E-5   -8.928093E-6   8.928093E-6   8.042445E-5   8.091850E-5   -6.334592E+0   8.366541E+1   
5.603050E+2   5.003661E+1   5.003661E+1   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   6.683510E-2   -6.254494E-2   8.205544E-5   -8.543199E-6   8.543199E-6   8.205544E-5   8.249898E-5   -5.943932E+0   8.405607E+1   
5.825840E+2   5.002200E+1   5.002200E+1   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   6.776408E-2   -6.514286E-2   8.432178E-5   -7.531857E-6   7.531857E-6   8.432178E-5   8.465750E-5   -5.104273E+0   8.489573E+1   
6.048780E+2   5.002300E+1   5.002300E+1   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   6.961711E-2   -6.538307E-2   8.562385E-5   -8.745375E-6   8.745375E-6   8.562385E-5   8.606931E-5   -5.831804E+0   8.416820E+1   
6.271280E+2   5.004449E+1   5.004449E+1   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   7.073291E-2   -6.699649E-2   8.736450E-5   -8.515843E-6   8.515843E-6   8.736450E-5   8.777856E-5   -5.567311E+0   8.443269E+1   
6.494100E+2   5.003869E+1   5.003869E+1   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   7.281205E-2   -6.911950E-2   9.003262E-5   -8.665680E-6   8.665680E-6   9.003262E-5   9.044869E-5   -5.497809E+0   8.450219E+1   
6.716120E+2   5.004531E+1   5.004531E+1   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   7.291728E-2   -7.098264E-2   9.131111E-5   -7.525439E-6   7.525439E-6   9.131111E-5   9.162069E-5   -4.711405E+0   8.528860E+1   
6.941860E+2   5.003961E+1   5.003961E+1   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   7.454511E-2   -7.323329E-2   9.378334E-5   -7.258021E-6   7.258021E-6   9.378334E-5   9.406377E-5   -4.425378E+0   8.557462E+1   
7.164580E+2   5.004519E+1   5.004519E+1   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   7.332194E-2   -7.476694E-2   9.402597E-5   -5.350672E-6   5.350672E-6   9.402597E-5   9.417809E-5   -3.256979E+0   8.674302E+1   
7.384520E+2   5.002981E+1   5.002981E+1   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   7.398092E-2   -7.557440E-2   9.495927E-5   -5.310179E-6   5.310179E-6   9.495927E-5   9.510763E-5   -3.200680E+0   8.679932E+1   
7.606330E+2   5.005410E+1   5.005410E+1   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   7.664849E-2   -7.677734E-2   9.739195E-5   -6.496748E-6   6.496748E-6   9.739195E-5   9.760840E-5   -3.816389E+0   8.618361E+1   
7.828260E+2   5.001739E+1   5.001739E+1   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   7.877764E-2   -7.955474E-2   1.005172E-4   -6.255744E-6   6.255744E-6   1.005172E-4   1.007117E-4   -3.561243E+0   8.643876E+1   
8.050950E+2   5.003350E+1   5.003350E+1   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   8.045027E-2   -8.062851E-2   1.022506E-4   -6.790874E-6   6.790874E-6   1.022506E-4   1.024759E-4   -3.799663E+0   8.620034E+1   
8.273640E+2   5.001110E+1   5.001110E+1   1.148000E+3   1.148000E+3   9.000000E+1   1.149000E+3   1.149000E+3   8.094696E-2   -8.220542E-2   1.035847E-4   -6.127309E-6   6.127309E-6   1.035847E-4   1.037658E-4   -3.385252E+0   8.661475E+1   
8.496710E+2   5.001699E+1   5.001699E+1   1.098000E+3   1.098000E+3   9.000000E+1   1.099000E+3   1.099000E+3   8.142002E-2   -8.444502E-2   1.053358E-4   -5.013010E-6   5.013010E-6   1.053358E-4   1.054550E-4   -2.724693E+0   8.727531E+1   
8.719700E+2   5.001141E+1   5.001141E+1   1.048000E+3   1.048000E+3   9.000000E+1   1.049000E+3   1.049000E+3   8.328750E-2   -8.552063E-2   1.071909E-4   -5.691050E-6   5.691050E-6   1.071909E-4   1.073419E-4   -3.039132E+0   8.696087E+1   
8.941020E+2   5.003100E+1   5.003100E+1   9.980000E+2   9.980000E+2   9.000000E+1   9.990000E+2   9.990000E+2   8.402471E-2   -8.798570E-2   1.092522E-4   -4.624718E-6   4.624718E-6   1.092522E-4   1.093500E-4   -2.423922E+0   8.757608E+1   
9.159460E+2   5.000030E+1   5.000030E+1   9.480000E+2   9.480000E+2   9.000000E+1   9.480000E+2   9.480000E+2   8.528806E-2   -8.901929E-2   1.107064E-4   -4.883398E-6   4.883398E-6   1.107064E-4   1.108140E-4   -2.525751E+0   8.747425E+1   
9.377750E+2   5.000271E+1   5.000271E+1   8.980000E+2   8.980000E+2   9.000000E+1   8.990000E+2   8.990000E+2   8.534145E-2   -9.162646E-2   1.124374E-4   -3.218394E-6   3.218394E-6   1.124374E-4   1.124835E-4   -1.639579E+0   8.836042E+1   
9.595890E+2   5.001150E+1   5.001150E+1   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   8.780563E-2   -9.227750E-2   1.143849E-4   -4.615350E-6   4.615350E-6   1.143849E-4   1.144780E-4   -2.310591E+0   8.768941E+1   
9.814360E+2   5.003411E+1   5.003411E+1   7.980000E+2   7.980000E+2   9.000000E+1   7.990000E+2   7.990000E+2   8.813420E-2   -9.443500E-2   1.159932E-4   -3.447860E-6   3.447860E-6   1.159932E-4   1.160444E-4   -1.702597E+0   8.829740E+1   
1.003324E+3   5.003649E+1   5.003649E+1   7.480000E+2   7.480000E+2   9.000000E+1   7.480000E+2   7.480000E+2   8.970744E-2   -9.515784E-2   1.174366E-4   -4.138898E-6   4.138898E-6   1.174366E-4   1.175095E-4   -2.018478E+0   8.798152E+1   
1.025206E+3   5.003411E+1   5.003411E+1   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   9.084168E-2   -9.742572E-2   1.196149E-4   -3.495144E-6   3.495144E-6   1.196149E-4   1.196660E-4   -1.673705E+0   8.832630E+1   
1.047025E+3   5.001479E+1   5.001479E+1   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   9.235451E-2   -9.756228E-2   1.206392E-4   -4.524804E-6   4.524804E-6   1.206392E-4   1.207240E-4   -2.147982E+0   8.785202E+1   
1.068895E+3   5.002429E+1   5.002429E+1   5.980000E+2   5.980000E+2   9.000000E+1   5.990000E+2   5.990000E+2   9.249657E-2   -9.913703E-2   1.217526E-4   -3.600345E-6   3.600345E-6   1.217526E-4   1.218058E-4   -1.693799E+0   8.830620E+1   
1.090825E+3   5.001751E+1   5.001751E+1   5.480000E+2   5.480000E+2   9.000000E+1   5.480000E+2   5.480000E+2   9.328013E-2   -1.028532E-1   1.246574E-4   -1.750342E-6   1.750342E-6   1.246574E-4   1.246696E-4   -8.044500E-1   8.919555E+1   
1.112669E+3   5.000219E+1   5.000219E+1   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   9.379065E-2   -1.037245E-1   1.255404E-4   -1.558322E-6   1.558322E-6   1.255404E-4   1.255501E-4   -7.111709E-1   8.928883E+1   
1.134747E+3   5.003781E+1   5.003781E+1   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   9.420303E-2   -1.051944E-1   1.267527E-4   -9.023732E-7   9.023732E-7   1.267527E-4   1.267559E-4   -4.078911E-1   8.959211E+1   
1.156541E+3   5.002581E+1   5.002581E+1   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   9.625223E-2   -1.074662E-1   1.294992E-4   -9.327950E-7   9.327950E-7   1.294992E-4   1.295026E-4   -4.126998E-1   8.958730E+1   
1.178403E+3   5.003311E+1   5.003311E+1   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   9.720143E-2   -1.082476E-1   1.305950E-4   -1.124001E-6   1.124001E-6   1.305950E-4   1.305998E-4   -4.931196E-1   8.950688E+1   
1.200215E+3   5.002889E+1   5.002889E+1   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   9.731311E-2   -1.088575E-1   1.310612E-4   -8.078513E-7   8.078513E-7   1.310612E-4   1.310637E-4   -3.531623E-1   8.964684E+1   
1.222094E+3   5.003079E+1   5.003079E+1   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   1.001605E-1   -1.095708E-1   1.332862E-4   -2.447535E-6   2.447535E-6   1.332862E-4   1.333086E-4   -1.052005E+0   8.894800E+1   
1.243947E+3   5.002160E+1   5.002160E+1   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   1.010812E-1   -1.121938E-1   1.355638E-4   -1.413619E-6   1.413619E-6   1.355638E-4   1.355711E-4   -5.974419E-1   8.940256E+1   
1.265793E+3   5.004449E+1   5.004449E+1   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   1.004148E-1   -1.144638E-1   1.366302E-4   5.632536E-7   -5.632536E-7   1.366302E-4   1.366314E-4   2.361987E-1   9.023620E+1   
1.287663E+3   5.000851E+1   5.000851E+1   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   1.016721E-1   -1.153885E-1   1.380097E-4   2.378970E-7   -2.378970E-7   1.380097E-4   1.380099E-4   9.876463E-2   9.009876E+1   
1.309395E+3   5.001299E+1   5.001299E+1   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   1.027624E-1   -1.167565E-1   1.395748E-4   3.257902E-7   -3.257902E-7   1.395748E-4   1.395752E-4   1.337374E-1   9.013374E+1   
1.342530E+3   5.002361E+1   5.002361E+1   4.700000E+1   4.700000E+1   9.000000E+1   4.700000E+1   4.700000E+1   1.038445E-1   -1.170556E-1   1.404386E-4   -2.789638E-7   2.789638E-7   1.404386E-4   1.404388E-4   -1.138108E-1   8.988619E+1   
1.363958E+3   5.004739E+1   5.004739E+1   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   1.033677E-1   -1.177575E-1   1.406010E-4   5.325585E-7   -5.325585E-7   1.406010E-4   1.406020E-4   2.170199E-1   9.021702E+1   
1.382936E+3   5.003680E+1   5.003680E+1   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   1.040807E-1   -1.173682E-1   1.407882E-4   -2.493089E-7   2.493089E-7   1.407882E-4   1.407884E-4   -1.014597E-1   8.989854E+1   
1.405362E+3   5.001849E+1   5.001849E+1   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   1.032401E-1   -1.175216E-1   1.403684E-4   4.727194E-7   -4.727194E-7   1.403684E-4   1.403692E-4   1.929545E-1   9.019295E+1   
1.424470E+3   5.002480E+1   5.002480E+1   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   1.035601E-1   -1.162960E-1   1.397680E-4   -5.652445E-7   5.652445E-7   1.397680E-4   1.397692E-4   -2.317122E-1   8.976829E+1   
1.446909E+3   5.003411E+1   5.003411E+1   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   1.037426E-1   -1.173992E-1   1.405994E-4   2.101698E-8   -2.101698E-8   1.405994E-4   1.405994E-4   8.564650E-3   9.000856E+1   
1.465967E+3   5.003900E+1   5.003900E+1   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   1.035024E-1   -1.176762E-1   1.406313E-4   3.798035E-7   -3.798035E-7   1.406313E-4   1.406318E-4   1.547385E-1   9.015474E+1   
1.488398E+3   5.002261E+1   5.002261E+1   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   1.031695E-1   -1.178606E-1   1.405456E-4   7.465494E-7   -7.465494E-7   1.405456E-4   1.405476E-4   3.043406E-1   9.030434E+1   
1.507413E+3   5.003231E+1   5.003231E+1   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   1.036668E-1   -1.177247E-1   1.407645E-4   2.898705E-7   -2.898705E-7   1.407645E-4   1.407648E-4   1.179866E-1   9.011799E+1   
1.529852E+3   5.005721E+1   5.005721E+1   2.900000E+1   2.900000E+1   9.000000E+1   2.900000E+1   2.900000E+1   1.028603E-1   -1.178222E-1   1.403294E-4   9.501931E-7   -9.501931E-7   1.403294E-4   1.403326E-4   3.879530E-1   9.038795E+1   
1.551270E+3   5.003909E+1   5.003909E+1   2.700000E+1   2.700000E+1   9.000000E+1   2.700000E+1   2.700000E+1   1.036303E-1   -1.179548E-1   1.408918E-4   4.672943E-7   -4.672943E-7   1.408918E-4   1.408926E-4   1.900316E-1   9.019003E+1   
1.572615E+3   5.003259E+1   5.003259E+1   2.500000E+1   2.500000E+1   9.000000E+1   2.500000E+1   2.500000E+1   1.036217E-1   -1.175247E-1   1.406064E-4   1.924496E-7   -1.924496E-7   1.406064E-4   1.406065E-4   7.842135E-2   9.007842E+1   
1.593977E+3   5.004031E+1   5.004031E+1   2.200000E+1   2.200000E+1   9.000000E+1   2.400000E+1   2.400000E+1   1.042636E-1   -1.189181E-1   1.419107E-4   6.287445E-7   -6.287445E-7   1.419107E-4   1.419121E-4   2.538509E-1   9.025385E+1   
1.612959E+3   5.002569E+1   5.002569E+1   2.300000E+1   2.300000E+1   9.000000E+1   2.300000E+1   2.300000E+1   1.041654E-1   -1.184300E-1   1.415321E-4   3.822575E-7   -3.822575E-7   1.415321E-4   1.415326E-4   1.547471E-1   9.015475E+1   
1.635011E+3   5.001739E+1   5.001739E+1   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   1.036711E-1   -1.183416E-1   1.411690E-4   6.900369E-7   -6.900369E-7   1.411690E-4   1.411707E-4   2.800607E-1   9.028006E+1   
1.653988E+3   5.002789E+1   5.002789E+1   1.900000E+1   1.900000E+1   9.000000E+1   2.000000E+1   2.000000E+1   1.041605E-1   -1.172829E-1   1.407820E-4   -3.640669E-7   3.640669E-7   1.407820E-4   1.407825E-4   -1.481685E-1   8.985183E+1   
1.676058E+3   5.002160E+1   5.002160E+1   1.500000E+1   1.500000E+1   9.000000E+1   1.600000E+1   1.600000E+1   1.046102E-1   -1.188086E-1   1.420537E-4   3.007330E-7   -3.007330E-7   1.420537E-4   1.420540E-4   1.212971E-1   9.012130E+1   
1.697430E+3   5.000479E+1   5.000479E+1   1.300000E+1   1.300000E+1   9.000000E+1   1.300000E+1   1.300000E+1   1.038356E-1   -1.175326E-1   1.407438E-4   3.950265E-8   -3.950265E-8   1.407438E-4   1.407438E-4   1.608124E-2   9.001608E+1   
1.718796E+3   5.001470E+1   5.001470E+1   1.100000E+1   1.100000E+1   9.000000E+1   1.100000E+1   1.100000E+1   1.031140E-1   -1.186945E-1   1.410543E-4   1.332782E-6   -1.332782E-6   1.410543E-4   1.410606E-4   5.413551E-1   9.054136E+1   
1.739928E+3   5.000121E+1   5.000121E+1   9.000000E+0   9.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   1.047670E-1   -1.183938E-1   1.418805E-4   -8.639189E-8   8.639189E-8   1.418805E-4   1.418805E-4   -3.488774E-2   8.996511E+1   
1.760960E+3   5.001309E+1   5.001309E+1   7.000000E+0   7.000000E+0   9.000000E+1   7.000000E+0   7.000000E+0   1.049630E-1   -1.174633E-1   1.413957E-4   -8.397400E-7   8.397400E-7   1.413957E-4   1.413982E-4   -3.402720E-1   8.965973E+1   
1.782048E+3   5.002279E+1   5.002279E+1   5.000000E+0   5.000000E+0   9.000000E+1   6.000000E+0   6.000000E+0   1.050207E-1   -1.181680E-1   1.418903E-4   -4.216705E-7   4.216705E-7   1.418903E-4   1.418909E-4   -1.702714E-1   8.982973E+1   
1.803053E+3   4.999749E+1   4.999749E+1   3.000000E+0   3.000000E+0   9.000000E+1   3.000000E+0   3.000000E+0   1.052474E-1   -1.181180E-1   1.419979E-4   -6.220688E-7   6.220688E-7   1.419979E-4   1.419993E-4   -2.510015E-1   8.974900E+1   
1.824049E+3   5.001919E+1   5.001919E+1   1.000000E+0   1.000000E+0   9.000000E+1   2.000000E+0   2.000000E+0   1.027069E-1   -1.194314E-1   1.412826E-4   2.115659E-6   -2.115659E-6   1.412826E-4   1.412984E-4   8.579209E-1   9.085792E+1   
1.845071E+3   5.003600E+1   5.003600E+1   0.000000E+0   0.000000E+0   9.000000E+1   0.000000E+0   0.000000E+0   1.052140E-1   -1.183404E-1   1.421221E-4   -4.519067E-7   4.519067E-7   1.421221E-4   1.421228E-4   -1.821833E-1   8.981782E+1   
1.867124E+3   5.003631E+1   5.003631E+1   -1.000000E+0   -1.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   1.039147E-1   -1.187662E-1   1.415961E-4   7.874500E-7   -7.874500E-7   1.415961E-4   1.415983E-4   3.186322E-1   9.031863E+1   
1.888862E+3   5.000430E+1   5.000430E+1   -3.000000E+0   -3.000000E+0   9.000000E+1   -2.000000E+0   -2.000000E+0   1.046538E-1   -1.183693E-1   1.417945E-4   -1.872817E-8   1.872817E-8   1.417945E-4   1.417945E-4   -7.567604E-3   8.999243E+1   
1.910560E+3   5.005840E+1   5.005840E+1   -5.000000E+0   -5.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   1.059297E-1   -1.191464E-1   1.430895E-4   -4.544078E-7   4.544078E-7   1.430895E-4   1.430902E-4   -1.819530E-1   8.981805E+1   
1.932314E+3   5.002941E+1   5.002941E+1   -7.000000E+0   -7.000000E+0   9.000000E+1   -6.000000E+0   -6.000000E+0   1.050124E-1   -1.183732E-1   1.420188E-4   -2.813703E-7   2.813703E-7   1.420188E-4   1.420191E-4   -1.135153E-1   8.988648E+1   
1.954045E+3   5.003039E+1   5.003039E+1   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   1.042795E-1   -1.192442E-1   1.421330E-4   8.301530E-7   -8.301530E-7   1.421330E-4   1.421354E-4   3.346424E-1   9.033464E+1   
1.976287E+3   5.001830E+1   5.001830E+1   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   1.042571E-1   -1.192108E-1   1.420974E-4   8.248524E-7   -8.248524E-7   1.420974E-4   1.420997E-4   3.325891E-1   9.033259E+1   
1.998552E+3   5.003381E+1   5.003381E+1   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   1.039540E-1   -1.198026E-1   1.422954E-4   1.435957E-6   -1.435957E-6   1.422954E-4   1.423026E-4   5.781738E-1   9.057817E+1   
2.020770E+3   5.000631E+1   5.000631E+1   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   1.052634E-1   -1.187073E-1   1.423916E-4   -2.485650E-7   2.485650E-7   1.423916E-4   1.423918E-4   -1.000179E-1   8.989998E+1   
2.042953E+3   5.002429E+1   5.002429E+1   -1.700000E+1   -1.700000E+1   9.000000E+1   -1.600000E+1   -1.600000E+1   1.051928E-1   -1.186714E-1   1.423246E-4   -2.198438E-7   2.198438E-7   1.423246E-4   1.423248E-4   -8.850270E-2   8.991150E+1   
2.064847E+3   5.001541E+1   5.001541E+1   -1.900000E+1   -1.900000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   1.040325E-1   -1.187396E-1   1.416516E-4   6.828865E-7   -6.828865E-7   1.416516E-4   1.416532E-4   2.762144E-1   9.027621E+1   
2.086732E+3   5.003820E+1   5.003820E+1   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   1.047983E-1   -1.185582E-1   1.420069E-4   -2.045063E-9   2.045063E-9   1.420069E-4   1.420069E-4   -8.251249E-4   8.999917E+1   
2.108927E+3   5.003240E+1   5.003240E+1   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   1.058905E-1   -1.190292E-1   1.429889E-4   -5.019790E-7   5.019790E-7   1.429889E-4   1.429898E-4   -2.011426E-1   8.979886E+1   
2.131201E+3   4.999691E+1   4.999691E+1   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   1.051327E-1   -1.196909E-1   1.429514E-4   4.911368E-7   -4.911368E-7   1.429514E-4   1.429522E-4   1.968498E-1   9.019685E+1   
2.153432E+3   5.000891E+1   5.000891E+1   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   1.052793E-1   -1.195231E-1   1.429327E-4   2.729583E-7   -2.729583E-7   1.429327E-4   1.429330E-4   1.094175E-1   9.010942E+1   
2.175663E+3   5.001431E+1   5.001431E+1   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   1.052760E-1   -1.203076E-1   1.434416E-4   7.883202E-7   -7.883202E-7   1.434416E-4   1.434437E-4   3.148806E-1   9.031488E+1   
2.197903E+3   5.001980E+1   5.001980E+1   -3.100000E+1   -3.100000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   1.044314E-1   -1.188196E-1   1.419503E-4   4.402311E-7   -4.402311E-7   1.419503E-4   1.419510E-4   1.776911E-1   9.017769E+1   
2.219822E+3   5.002480E+1   5.002480E+1   -3.300000E+1   -3.300000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   1.056380E-1   -1.188936E-1   1.427445E-4   -4.038809E-7   4.038809E-7   1.427445E-4   1.427450E-4   -1.621121E-1   8.983789E+1   
2.241700E+3   5.001000E+1   5.001000E+1   -3.500000E+1   -3.500000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   1.055187E-1   -1.196342E-1   1.431530E-4   1.685747E-7   -1.685747E-7   1.431530E-4   1.431531E-4   6.747056E-2   9.006747E+1   
2.263580E+3   5.002471E+1   5.002471E+1   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   1.048900E-1   -1.201695E-1   1.431131E-4   9.835109E-7   -9.835109E-7   1.431131E-4   1.431164E-4   3.937456E-1   9.039375E+1   
2.285823E+3   5.001629E+1   5.001629E+1   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   1.058337E-1   -1.198907E-1   1.435149E-4   1.032454E-7   -1.032454E-7   1.435149E-4   1.435149E-4   4.121890E-2   9.004122E+1   
2.308135E+3   5.001931E+1   5.001931E+1   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   1.052069E-1   -1.202849E-1   1.433841E-4   8.245268E-7   -8.245268E-7   1.433841E-4   1.433865E-4   3.294743E-1   9.032947E+1   
2.330374E+3   5.002950E+1   5.002950E+1   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   1.055297E-1   -1.202652E-1   1.435709E-4   5.729851E-7   -5.729851E-7   1.435709E-4   1.435720E-4   2.286638E-1   9.022866E+1   
2.352628E+3   5.001739E+1   5.001739E+1   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   1.051367E-1   -1.202717E-1   1.433321E-4   8.678731E-7   -8.678731E-7   1.433321E-4   1.433347E-4   3.469206E-1   9.034692E+1   
2.374849E+3   5.001422E+1   5.001422E+1   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   1.058791E-1   -1.206533E-1   1.440397E-4   5.682606E-7   -5.682606E-7   1.440397E-4   1.440408E-4   2.260403E-1   9.022604E+1   
2.397032E+3   5.001769E+1   5.001769E+1   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   1.055877E-1   -1.198983E-1   1.433677E-4   2.902104E-7   -2.902104E-7   1.433677E-4   1.433680E-4   1.159801E-1   9.011598E+1   
2.430398E+3   5.001730E+1   5.001730E+1   -9.900000E+1   -9.900000E+1   9.000000E+1   -9.900000E+1   -9.900000E+1   1.071680E-1   -1.208503E-1   1.449648E-4   -2.562423E-7   2.562423E-7   1.449648E-4   1.449650E-4   -1.012769E-1   8.989872E+1   
2.452521E+3   5.003411E+1   5.003411E+1   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   1.076346E-1   -1.236323E-1   1.470651E-4   1.217403E-6   -1.217403E-6   1.470651E-4   1.470702E-4   4.742827E-1   9.047428E+1   
2.474227E+3   5.001589E+1   5.001589E+1   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   1.089001E-1   -1.250055E-1   1.487419E-4   1.179152E-6   -1.179152E-6   1.487419E-4   1.487466E-4   4.542029E-1   9.045420E+1   
2.495949E+3   5.001019E+1   5.001019E+1   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   1.097603E-1   -1.269217E-1   1.505217E-4   1.795661E-6   -1.795661E-6   1.505217E-4   1.505325E-4   6.834821E-1   9.068348E+1   
2.518125E+3   5.004171E+1   5.004171E+1   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   1.115790E-1   -1.272061E-1   1.518314E-4   6.364449E-7   -6.364449E-7   1.518314E-4   1.518327E-4   2.401704E-1   9.024017E+1   
2.539817E+3   5.003060E+1   5.003060E+1   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   1.118033E-1   -1.289165E-1   1.530840E-4   1.588756E-6   -1.588756E-6   1.530840E-4   1.530922E-4   5.946130E-1   9.059461E+1   
2.561429E+3   5.002630E+1   5.002630E+1   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   1.119100E-1   -1.305127E-1   1.541896E-4   2.553374E-6   -2.553374E-6   1.541896E-4   1.542107E-4   9.487293E-1   9.094873E+1   
2.583605E+3   5.002429E+1   5.002429E+1   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   1.151645E-1   -1.315246E-1   1.568606E-4   8.077959E-7   -8.077959E-7   1.568606E-4   1.568627E-4   2.950574E-1   9.029506E+1   
2.605288E+3   4.999700E+1   4.999700E+1   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   1.144883E-1   -1.329290E-1   1.573573E-4   2.226105E-6   -2.226105E-6   1.573573E-4   1.573730E-4   8.104991E-1   9.081050E+1   
2.626984E+3   5.000140E+1   5.000140E+1   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   1.164665E-1   -1.343440E-1   1.595019E-4   1.688020E-6   -1.688020E-6   1.595019E-4   1.595108E-4   6.063428E-1   9.060634E+1   
2.649367E+3   5.000549E+1   5.000549E+1   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   1.162202E-1   -1.355950E-1   1.601644E-4   2.688148E-6   -2.688148E-6   1.601644E-4   1.601869E-4   9.615439E-1   9.096154E+1   
2.671060E+3   5.001699E+1   5.001699E+1   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.490000E+2   -6.490000E+2   1.169200E-1   -1.374066E-1   1.617769E-4   3.354938E-6   -3.354938E-6   1.617769E-4   1.618117E-4   1.188033E+0   9.118803E+1   
2.692725E+3   5.001431E+1   5.001431E+1   -7.000000E+2   -7.000000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   1.173903E-1   -1.390388E-1   1.631307E-4   4.074136E-6   -4.074136E-6   1.631307E-4   1.631815E-4   1.430647E+0   9.143065E+1   
2.714375E+3   5.001660E+1   5.001660E+1   -7.510000E+2   -7.510000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   1.203036E-1   -1.414796E-1   1.665215E-4   3.515115E-6   -3.515115E-6   1.665215E-4   1.665586E-4   1.209281E+0   9.120928E+1   
2.736106E+3   5.000121E+1   5.000121E+1   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   1.197228E-1   -1.422040E-1   1.666342E-4   4.418203E-6   -4.418203E-6   1.666342E-4   1.666928E-4   1.518806E+0   9.151881E+1   
2.757839E+3   5.003689E+1   5.003689E+1   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.490000E+2   -8.490000E+2   1.200112E-1   -1.433713E-1   1.675728E-4   4.968094E-6   -4.968094E-6   1.675728E-4   1.676464E-4   1.698172E+0   9.169817E+1   
2.779570E+3   5.004171E+1   5.004171E+1   -9.000000E+2   -9.000000E+2   9.000000E+1   -8.990000E+2   -8.990000E+2   1.220633E-1   -1.440901E-1   1.693096E-4   3.920216E-6   -3.920216E-6   1.693096E-4   1.693550E-4   1.326396E+0   9.132640E+1   
2.801305E+3   5.000381E+1   5.000381E+1   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   1.233445E-1   -1.468319E-1   1.718874E-4   4.765134E-6   -4.765134E-6   1.718874E-4   1.719535E-4   1.587971E+0   9.158797E+1   
2.823008E+3   5.000189E+1   5.000189E+1   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   1.241719E-1   -1.482613E-1   1.733299E-4   5.087633E-6   -5.087633E-6   1.733299E-4   1.734046E-4   1.681281E+0   9.168128E+1   
2.845521E+3   5.001650E+1   5.001650E+1   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   1.235663E-1   -1.502223E-1   1.742327E-4   6.817604E-6   -6.817604E-6   1.742327E-4   1.743660E-4   2.240801E+0   9.224080E+1   
2.867314E+3   5.001989E+1   5.001989E+1   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   1.269226E-1   -1.510816E-1   1.768674E-4   4.896977E-6   -4.896977E-6   1.768674E-4   1.769352E-4   1.585959E+0   9.158596E+1   
2.889197E+3   5.004861E+1   5.004861E+1   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   1.263229E-1   -1.512136E-1   1.765825E-4   5.426856E-6   -5.426856E-6   1.765825E-4   1.766659E-4   1.760300E+0   9.176030E+1   
2.911577E+3   5.001650E+1   5.001650E+1   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   1.265527E-1   -1.542075E-1   1.786745E-4   7.214257E-6   -7.214257E-6   1.786745E-4   1.788201E-4   2.312149E+0   9.231215E+1   
2.933455E+3   5.002319E+1   5.002319E+1   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   1.275083E-1   -1.546950E-1   1.795828E-4   6.826154E-6   -6.826154E-6   1.795828E-4   1.797125E-4   2.176832E+0   9.217683E+1   
2.955567E+3   5.004220E+1   5.004220E+1   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   1.307695E-1   -1.558111E-1   1.823260E-4   5.143721E-6   -5.143721E-6   1.823260E-4   1.823985E-4   1.615981E+0   9.161598E+1   
2.977921E+3   5.000451E+1   5.000451E+1   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   1.298347E-1   -1.581281E-1   1.832570E-4   7.349862E-6   -7.349862E-6   1.832570E-4   1.834044E-4   2.296722E+0   9.229672E+1   
2.999962E+3   5.000289E+1   5.000289E+1   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   1.311183E-1   -1.587576E-1   1.844606E-4   6.812029E-6   -6.812029E-6   1.844606E-4   1.845864E-4   2.114940E+0   9.211494E+1   
3.021736E+3   5.002780E+1   5.002780E+1   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   1.325980E-1   -1.609607E-1   1.868103E-4   7.157936E-6   -7.157936E-6   1.868103E-4   1.869473E-4   2.194307E+0   9.219431E+1   
3.044103E+3   5.004659E+1   5.004659E+1   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   1.327486E-1   -1.622204E-1   1.877238E-4   7.870083E-6   -7.870083E-6   1.877238E-4   1.878887E-4   2.400647E+0   9.240065E+1   
3.066195E+3   5.001510E+1   5.001510E+1   -1.550000E+3   -1.550000E+3   9.000000E+1   -1.548000E+3   -1.548000E+3   1.340089E-1   -1.636279E-1   1.894197E-4   7.858146E-6   -7.858146E-6   1.894197E-4   1.895826E-4   2.375574E+0   9.237557E+1   
3.088318E+3   5.002941E+1   5.002941E+1   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   1.347857E-1   -1.649082E-1   1.907338E-4   8.120571E-6   -8.120571E-6   1.907338E-4   1.909066E-4   2.437920E+0   9.243792E+1   
3.111169E+3   5.002319E+1   5.002319E+1   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.648000E+3   -1.648000E+3   1.348606E-1   -1.665253E-1   1.918333E-4   9.122440E-6   -9.122440E-6   1.918333E-4   1.920500E-4   2.722593E+0   9.272259E+1   
3.133534E+3   5.002191E+1   5.002191E+1   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.698000E+3   -1.698000E+3   1.372336E-1   -1.687916E-1   1.947764E-4   8.848890E-6   -8.848890E-6   1.947764E-4   1.949773E-4   2.601217E+0   9.260122E+1   
3.155661E+3   4.998800E+1   4.998800E+1   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.748000E+3   -1.748000E+3   1.389145E-1   -1.697714E-1   1.964538E-4   8.246259E-6   -8.246259E-6   1.964538E-4   1.966268E-4   2.403612E+0   9.240361E+1   
3.178968E+3   5.002639E+1   5.002639E+1   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.798000E+3   -1.798000E+3   1.387538E-1   -1.714223E-1   1.974296E-4   9.444429E-6   -9.444429E-6   1.974296E-4   1.976554E-4   2.738767E+0   9.273877E+1   
3.201335E+3   5.001620E+1   5.001620E+1   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.848000E+3   -1.848000E+3   1.391790E-1   -1.726669E-1   1.985031E-4   9.943641E-6   -9.943641E-6   1.985031E-4   1.987520E-4   2.867727E+0   9.286773E+1   
3.223370E+3   5.003109E+1   5.003109E+1   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   1.405317E-1   -1.746860E-1   2.006544E-4   1.026316E-5   -1.026316E-5   2.006544E-4   2.009167E-4   2.928039E+0   9.292804E+1   
3.246505E+3   5.002310E+1   5.002310E+1   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.948000E+3   -1.948000E+3   1.426096E-1   -1.766801E-1   2.032378E-4   1.003001E-5   -1.003001E-5   2.032378E-4   2.034851E-4   2.825317E+0   9.282532E+1   
3.268827E+3   5.003579E+1   5.003579E+1   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   1.434812E-1   -1.770173E-1   2.039962E-4   9.605755E-6   -9.605755E-6   2.039962E-4   2.042223E-4   2.695947E+0   9.269595E+1   
3.306403E+3   5.000359E+1   5.000359E+1   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.525429E-1   -1.949031E-1   2.212474E-4   1.459665E-5   -1.459665E-5   2.212474E-4   2.217284E-4   3.774581E+0   9.377458E+1   
3.332576E+3   5.002221E+1   5.002221E+1   -2.999000E+3   -2.999000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.629054E-1   -2.092383E-1   2.369904E-4   1.630416E-5   -1.630416E-5   2.369904E-4   2.375506E-4   3.935560E+0   9.393556E+1   
3.357762E+3   5.000701E+1   5.000701E+1   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.738377E-1   -2.281827E-1   2.560876E-4   2.060368E-5   -2.060368E-5   2.560876E-4   2.569151E-4   4.599858E+0   9.459986E+1   
3.383369E+3   5.004312E+1   5.004312E+1   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   1.815477E-1   -2.425470E-1   2.702096E-4   2.429211E-5   -2.429211E-5   2.702096E-4   2.712993E-4   5.137137E+0   9.513714E+1   
3.409519E+3   5.001891E+1   5.001891E+1   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   1.936513E-1   -2.574353E-1   2.873892E-4   2.507336E-5   -2.507336E-5   2.873892E-4   2.884809E-4   4.986164E+0   9.498616E+1   
3.434698E+3   5.003179E+1   5.003179E+1   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   1.975982E-1   -2.688530E-1   2.972656E-4   2.961870E-5   -2.961870E-5   2.972656E-4   2.987375E-4   5.690009E+0   9.569001E+1   
3.459836E+3   5.001211E+1   5.001211E+1   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   2.010589E-1   -2.769367E-1   3.046699E-4   3.234399E-5   -3.234399E-5   3.046699E-4   3.063819E-4   6.059866E+0   9.605987E+1   
3.485516E+3   5.004049E+1   5.004049E+1   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   1.931475E-1   -2.717506E-1   2.964011E-4   3.480495E-5   -3.480495E-5   2.964011E-4   2.984376E-4   6.697296E+0   9.669730E+1   
3.510827E+3   5.002831E+1   5.002831E+1   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.762408E-1   -2.535927E-1   2.741225E-4   3.543863E-5   -3.543863E-5   2.741225E-4   2.764038E-4   7.366354E+0   9.736635E+1   
3.535567E+3   5.001220E+1   5.001220E+1   -7.000000E+3   -7.000000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.581201E-1   -2.355561E-1   2.511724E-4   3.704944E-5   -3.704944E-5   2.511724E-4   2.538902E-4   8.390963E+0   9.839096E+1   
3.560783E+3   5.002761E+1   5.002761E+1   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.443166E-1   -2.211387E-1   2.332486E-4   3.783324E-5   -3.783324E-5   2.332486E-4   2.362969E-4   9.213217E+0   9.921322E+1   
3.586453E+3   5.002160E+1   5.002160E+1   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.347173E-1   -2.125252E-1   2.217040E-4   3.930189E-5   -3.930189E-5   2.217040E-4   2.251606E-4   1.005250E+1   1.000525E+2   
3.611678E+3   5.002120E+1   5.002120E+1   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.500000E+3   -8.500000E+3   1.277083E-1   -2.074999E-1   2.140978E-4   4.120056E-5   -4.120056E-5   2.140978E-4   2.180260E-4   1.089273E+1   1.008927E+2   
3.636879E+3   5.003051E+1   5.003051E+1   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.353880E-1   -2.193655E-1   2.265736E-4   4.327782E-5   -4.327782E-5   2.265736E-4   2.306698E-4   1.081381E+1   1.008138E+2   
3.662561E+3   5.004461E+1   5.004461E+1   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.343406E-1   -2.247242E-1   2.294161E-4   4.755588E-5   -4.755588E-5   2.294161E-4   2.342933E-4   1.171103E+1   1.017110E+2   
3.687761E+3   5.002151E+1   5.002151E+1   -9.999000E+3   -9.999000E+3   9.000000E+1   -9.999000E+3   -9.999000E+3   1.451170E-1   -2.396813E-1   2.458200E-4   4.936383E-5   -4.936383E-5   2.458200E-4   2.507275E-4   1.135471E+1   1.013547E+2   
3.724281E+3   5.005432E+1   5.005432E+1   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.323007E-1   -2.173759E-1   2.233691E-4   4.426052E-5   -4.426052E-5   2.233691E-4   2.277120E-4   1.120796E+1   1.012080E+2   
3.748463E+3   5.003341E+1   5.003341E+1   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.207892E-1   -2.013792E-1   2.058337E-4   4.231652E-5   -4.231652E-5   2.058337E-4   2.101385E-4   1.161734E+1   1.016173E+2   
3.773115E+3   5.003610E+1   5.003610E+1   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.093667E-1   -1.859703E-1   1.887361E-4   4.069110E-5   -4.069110E-5   1.887361E-4   1.930727E-4   1.216662E+1   1.021666E+2   
3.797767E+3   5.000921E+1   5.000921E+1   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.033030E-1   -1.710354E-1   1.752603E-4   3.541204E-5   -3.541204E-5   1.752603E-4   1.788021E-4   1.142305E+1   1.014230E+2   
3.822465E+3   4.998751E+1   4.998751E+1   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   8.903925E-2   -1.528748E-1   1.546140E-4   3.408905E-5   -3.408905E-5   1.546140E-4   1.583274E-4   1.243356E+1   1.024336E+2   
3.847604E+3   5.002859E+1   5.002859E+1   -7.000000E+3   -7.000000E+3   9.000000E+1   -6.999000E+3   -6.999000E+3   7.701665E-2   -1.353576E-1   1.357723E-4   3.152907E-5   -3.152907E-5   1.357723E-4   1.393850E-4   1.307352E+1   1.030735E+2   
3.872297E+3   5.001141E+1   5.001141E+1   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   6.507351E-2   -1.178882E-1   1.170108E-4   2.894160E-5   -2.894160E-5   1.170108E-4   1.205369E-4   1.389278E+1   1.038928E+2   
3.896494E+3   5.003140E+1   5.003140E+1   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   5.530095E-2   -1.038187E-1   1.018057E-4   2.697144E-5   -2.697144E-5   1.018057E-4   1.053179E-4   1.483852E+1   1.048385E+2   
3.921179E+3   5.002230E+1   5.002230E+1   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   4.231732E-2   -8.387132E-2   8.078705E-5   2.353349E-5   -2.353349E-5   8.078705E-5   8.414495E-5   1.624099E+1   1.062410E+2   
3.945837E+3   5.003869E+1   5.003869E+1   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   2.838126E-2   -6.446791E-2   5.953389E-5   2.115564E-5   -2.115564E-5   5.953389E-5   6.318105E-5   1.956290E+1   1.095629E+2   
3.970103E+3   5.001919E+1   5.001919E+1   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   2.059203E-2   -5.024712E-2   4.545637E-5   1.761965E-5   -1.761965E-5   4.545637E-5   4.875176E-5   2.118716E+1   1.111872E+2   
3.994826E+3   5.004330E+1   5.004330E+1   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   8.887828E-3   -3.381211E-2   2.751634E-5   1.553169E-5   -1.553169E-5   2.751634E-5   3.159719E-5   2.944270E+1   1.194427E+2   
4.019575E+3   5.001989E+1   5.001989E+1   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   -7.363094E-5   -1.905375E-2   1.236398E-5   1.251126E-5   -1.251126E-5   1.236398E-5   1.758977E-5   4.533923E+1   1.353392E+2   
4.043818E+3   4.999969E+1   4.999969E+1   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   -1.221808E-2   -1.918999E-3   -6.303967E-6   1.029146E-5   -1.029146E-5   -6.303967E-6   1.206873E-5   1.214893E+2   2.114893E+2   
4.068469E+3   5.000100E+1   5.000100E+1   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   -2.352684E-2   1.430827E-2   -2.386422E-5   8.046836E-6   -8.046836E-6   -2.386422E-5   2.518437E-5   1.613663E+2   2.513663E+2   
4.093075E+3   5.002410E+1   5.002410E+1   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.999000E+3   -1.999000E+3   -3.336786E-2   3.131943E-2   -4.102758E-5   4.204148E-6   -4.204148E-6   -4.102758E-5   4.124242E-5   1.741493E+2   2.641493E+2   
4.126774E+3   5.002450E+1   5.002450E+1   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.948000E+3   -1.948000E+3   -3.262787E-2   3.356974E-2   -4.203569E-5   2.185641E-6   -2.185641E-6   -4.203569E-5   4.209248E-5   1.770236E+2   2.670236E+2   
4.148804E+3   5.002621E+1   5.002621E+1   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.899000E+3   -1.899000E+3   -3.501165E-2   3.430911E-2   -4.399100E-5   3.465374E-6   -3.465374E-6   -4.399100E-5   4.412728E-5   1.754958E+2   2.654958E+2   
4.170935E+3   5.003201E+1   5.003201E+1   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.849000E+3   -1.849000E+3   -3.575287E-2   3.812438E-2   -4.693410E-5   1.519289E-6   -1.519289E-6   -4.693410E-5   4.695868E-5   1.781459E+2   2.681459E+2   
4.192754E+3   5.001360E+1   5.001360E+1   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.799000E+3   -1.799000E+3   -3.649348E-2   3.899321E-2   -4.795784E-5   1.499054E-6   -1.499054E-6   -4.795784E-5   4.798126E-5   1.782096E+2   2.682096E+2   
4.214789E+3   5.002499E+1   5.002499E+1   -1.750000E+3   -1.750000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   -3.682387E-2   4.026210E-2   -4.898852E-5   9.138523E-7   -9.138523E-7   -4.898852E-5   4.899704E-5   1.789313E+2   2.689313E+2   
4.236868E+3   5.000839E+1   5.000839E+1   -1.700000E+3   -1.700000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   -3.684351E-2   4.239001E-2   -5.038655E-5   -4.627882E-7   4.627882E-7   -5.038655E-5   5.038867E-5   -1.794738E+2   -8.947377E+1   
4.258710E+3   4.999929E+1   4.999929E+1   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   -3.808051E-2   4.285295E-2   -5.145282E-5   1.494771E-7   -1.494771E-7   -5.145282E-5   5.145304E-5   1.798335E+2   2.698335E+2   
4.280562E+3   5.002111E+1   5.002111E+1   -1.600000E+3   -1.600000E+3   9.000000E+1   -1.599000E+3   -1.599000E+3   -4.126839E-2   4.455018E-2   -5.452911E-5   1.397734E-6   -1.397734E-6   -5.452911E-5   5.454702E-5   1.785317E+2   2.685317E+2   
4.302554E+3   4.999941E+1   4.999941E+1   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   -4.009519E-2   4.624736E-2   -5.490914E-5   -5.795691E-7   5.795691E-7   -5.490914E-5   5.491220E-5   -1.793953E+2   -8.939526E+1   
4.324292E+3   4.999160E+1   4.999160E+1   -1.499000E+3   -1.499000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   -4.101190E-2   4.806089E-2   -5.665702E-5   -1.087171E-6   1.087171E-6   -5.665702E-5   5.666745E-5   -1.789007E+2   -8.890071E+1   
4.346355E+3   5.002099E+1   5.002099E+1   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   -4.195038E-2   4.909327E-2   -5.790961E-5   -1.067993E-6   1.067993E-6   -5.790961E-5   5.791946E-5   -1.789434E+2   -8.894345E+1   
4.368439E+3   5.002029E+1   5.002029E+1   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   -4.261644E-2   5.156145E-2   -5.992890E-5   -2.188980E-6   2.188980E-6   -5.992890E-5   5.996887E-5   -1.779081E+2   -8.790813E+1   
4.390343E+3   5.001711E+1   5.001711E+1   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   -4.389394E-2   5.154365E-2   -6.070712E-5   -1.232464E-6   1.232464E-6   -6.070712E-5   6.071963E-5   -1.788370E+2   -8.883695E+1   
4.412412E+3   5.001809E+1   5.001809E+1   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   -4.482874E-2   5.578598E-2   -6.404804E-5   -3.314569E-6   3.314569E-6   -6.404804E-5   6.413375E-5   -1.770375E+2   -8.703751E+1   
4.434451E+3   5.001620E+1   5.001620E+1   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   -4.661586E-2   5.503374E-2   -6.466300E-5   -1.500964E-6   1.500964E-6   -6.466300E-5   6.468042E-5   -1.786703E+2   -8.867028E+1   
4.456198E+3   4.999331E+1   4.999331E+1   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   -4.698799E-2   5.732363E-2   -6.638444E-5   -2.722787E-6   2.722787E-6   -6.638444E-5   6.644026E-5   -1.776513E+2   -8.765131E+1   
4.478298E+3   5.002551E+1   5.002551E+1   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   -4.892698E-2   5.862687E-2   -6.843200E-5   -2.140681E-6   2.140681E-6   -6.843200E-5   6.846548E-5   -1.782083E+2   -8.820827E+1   
4.500425E+3   5.002090E+1   5.002090E+1   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   -4.941631E-2   5.978380E-2   -6.948803E-5   -2.535117E-6   2.535117E-6   -6.948803E-5   6.953426E-5   -1.779106E+2   -8.791062E+1   
4.522546E+3   5.002889E+1   5.002889E+1   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   -4.958906E-2   6.170860E-2   -7.084843E-5   -3.665729E-6   3.665729E-6   -7.084843E-5   7.094320E-5   -1.770381E+2   -8.703813E+1   
4.544584E+3   5.001229E+1   5.001229E+1   -1.000000E+3   -1.000000E+3   9.000000E+1   -1.000000E+3   -1.000000E+3   -5.008883E-2   6.328736E-2   -7.218564E-5   -4.328238E-6   4.328238E-6   -7.218564E-5   7.231529E-5   -1.765687E+2   -8.656866E+1   
4.566479E+3   5.001721E+1   5.001721E+1   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   -5.120738E-2   6.461362E-2   -7.374096E-5   -4.367993E-6   4.367993E-6   -7.374096E-5   7.387022E-5   -1.766101E+2   -8.661009E+1   
4.588107E+3   5.001559E+1   5.001559E+1   -9.000000E+2   -9.000000E+2   9.000000E+1   -8.990000E+2   -8.990000E+2   -5.205446E-2   6.682682E-2   -7.570610E-5   -5.188395E-6   5.188395E-6   -7.570610E-5   7.588368E-5   -1.760795E+2   -8.607946E+1   
4.609975E+3   5.000240E+1   5.000240E+1   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   -5.372557E-2   6.711215E-2   -7.692509E-5   -4.138930E-6   4.138930E-6   -7.692509E-5   7.703636E-5   -1.769202E+2   -8.692019E+1   
4.631554E+3   5.000170E+1   5.000170E+1   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   -5.406335E-2   6.863720E-2   -7.812717E-5   -4.886133E-6   4.886133E-6   -7.812717E-5   7.827982E-5   -1.764213E+2   -8.642134E+1   
4.653188E+3   5.003579E+1   5.003579E+1   -7.500000E+2   -7.500000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   -5.529757E-2   7.039975E-2   -8.003816E-5   -5.125566E-6   5.125566E-6   -8.003816E-5   8.020211E-5   -1.763358E+2   -8.633584E+1   
4.675129E+3   5.000439E+1   5.000439E+1   -7.000000E+2   -7.000000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   -5.628822E-2   7.271203E-2   -8.215659E-5   -5.904552E-6   5.904552E-6   -8.215659E-5   8.236849E-5   -1.758892E+2   -8.588925E+1   
4.697029E+3   5.000439E+1   5.000439E+1   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.500000E+2   -6.500000E+2   -5.762736E-2   7.363118E-2   -8.358313E-5   -5.514998E-6   5.514998E-6   -8.358313E-5   8.376488E-5   -1.762250E+2   -8.622497E+1   
4.718650E+3   5.000329E+1   5.000329E+1   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   -5.776848E-2   7.543175E-2   -8.484308E-5   -6.587785E-6   6.587785E-6   -8.484308E-5   8.509845E-5   -1.755601E+2   -8.556008E+1   
4.740327E+3   5.003011E+1   5.003011E+1   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   -5.928249E-2   7.617971E-2   -8.626625E-5   -5.956971E-6   5.956971E-6   -8.626625E-5   8.647168E-5   -1.760498E+2   -8.604981E+1   
4.762268E+3   5.002130E+1   5.002130E+1   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   -5.961905E-2   7.771214E-2   -8.747238E-5   -6.709897E-6   6.709897E-6   -8.747238E-5   8.772935E-5   -1.756135E+2   -8.561350E+1   
4.783913E+3   4.999929E+1   4.999929E+1   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   -6.282288E-2   7.928199E-2   -9.047556E-5   -5.366574E-6   5.366574E-6   -9.047556E-5   9.063458E-5   -1.766055E+2   -8.660547E+1   
4.805534E+3   5.003011E+1   5.003011E+1   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   -6.226422E-2   8.120774E-2   -9.138439E-5   -7.038779E-6   7.038779E-6   -9.138439E-5   9.165507E-5   -1.755956E+2   -8.559555E+1   
4.827226E+3   5.001699E+1   5.001699E+1   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   -6.316957E-2   8.234377E-2   -9.268401E-5   -7.111858E-6   7.111858E-6   -9.268401E-5   9.295646E-5   -1.756122E+2   -8.561216E+1   
4.848903E+3   5.001849E+1   5.001849E+1   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   -6.437128E-2   8.467142E-2   -9.494293E-5   -7.744784E-6   7.744784E-6   -9.494293E-5   9.525829E-5   -1.753365E+2   -8.533653E+1   
4.870512E+3   5.000570E+1   5.000570E+1   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   -6.444828E-2   8.502699E-2   -9.522212E-5   -7.920292E-6   7.920292E-6   -9.522212E-5   9.555094E-5   -1.752453E+2   -8.524525E+1   
4.892126E+3   5.002520E+1   5.002520E+1   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   -6.550918E-2   8.686314E-2   -9.707388E-5   -8.336043E-6   8.336043E-6   -9.707388E-5   9.743115E-5   -1.750919E+2   -8.509187E+1   
4.913834E+3   5.002520E+1   5.002520E+1   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   -6.685783E-2   8.860419E-2   -9.904161E-5   -8.476790E-6   8.476790E-6   -9.904161E-5   9.940370E-5   -1.751081E+2   -8.510808E+1   
4.935452E+3   5.003399E+1   5.003399E+1   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   -6.817613E-2   8.925891E-2   -1.002831E-4   -7.929765E-6   7.929765E-6   -1.002831E-4   1.005961E-4   -1.754788E+2   -8.547881E+1   
4.956978E+3   5.000591E+1   5.000591E+1   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   -6.996625E-2   9.068028E-2   -1.023155E-4   -7.534994E-6   7.534994E-6   -1.023155E-4   1.025926E-4   -1.757881E+2   -8.578807E+1   
4.990016E+3   5.000561E+1   5.000561E+1   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   -6.742755E-2   9.103647E-2   -1.009780E-4   -9.645566E-6   9.645566E-6   -1.009780E-4   1.014376E-4   -1.745436E+2   -8.454358E+1   
5.012244E+3   5.002770E+1   5.002770E+1   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   -6.793866E-2   9.097664E-2   -1.012550E-4   -9.228413E-6   9.228413E-6   -1.012550E-4   1.016746E-4   -1.747924E+2   -8.479243E+1   
5.034510E+3   5.002349E+1   5.002349E+1   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   -6.871883E-2   9.118008E-2   -1.018698E-4   -8.784384E-6   8.784384E-6   -1.018698E-4   1.022479E-4   -1.750715E+2   -8.507149E+1   
5.056777E+3   5.002151E+1   5.002151E+1   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   -6.912595E-2   9.203971E-2   -1.026814E-4   -9.045264E-6   9.045264E-6   -1.026814E-4   1.030790E-4   -1.749658E+2   -8.496578E+1   
5.079031E+3   5.003619E+1   5.003619E+1   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   -6.945298E-2   9.162030E-2   -1.026104E-4   -8.529186E-6   8.529186E-6   -1.026104E-4   1.029643E-4   -1.752484E+2   -8.524838E+1   
5.101312E+3   5.003201E+1   5.003201E+1   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   -6.939993E-2   9.225328E-2   -1.029899E-4   -8.982245E-6   8.982245E-6   -1.029899E-4   1.033808E-4   -1.750156E+2   -8.501557E+1   
5.123548E+3   5.001721E+1   5.001721E+1   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   -6.852494E-2   9.201977E-2   -1.022968E-4   -9.476758E-6   9.476758E-6   -1.022968E-4   1.027348E-4   -1.747072E+2   -8.470724E+1   
5.145830E+3   5.001681E+1   5.001681E+1   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   -6.874767E-2   9.188109E-2   -1.023442E-4   -9.221349E-6   9.221349E-6   -1.023442E-4   1.027588E-4   -1.748515E+2   -8.485148E+1   
5.168121E+3   5.002029E+1   5.002029E+1   -3.100000E+1   -3.100000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   -6.885505E-2   9.169855E-2   -1.022917E-4   -9.022591E-6   9.022591E-6   -1.022917E-4   1.026889E-4   -1.749593E+2   -8.495930E+1   
5.189383E+3   5.003079E+1   5.003079E+1   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   -7.008774E-2   9.208450E-2   -1.033052E-4   -8.363178E-6   8.363178E-6   -1.033052E-4   1.036432E-4   -1.753717E+2   -8.537165E+1   
5.211570E+3   5.003799E+1   5.003799E+1   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   -6.893788E-2   9.200378E-2   -1.025417E-4   -9.160872E-6   9.160872E-6   -1.025417E-4   1.029501E-4   -1.748949E+2   -8.489486E+1   
5.233870E+3   5.001241E+1   5.001241E+1   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   -6.923578E-2   9.157703E-2   -1.024479E-4   -8.661542E-6   8.661542E-6   -1.024479E-4   1.028134E-4   -1.751674E+2   -8.516738E+1   
5.256142E+3   5.001461E+1   5.001461E+1   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   -6.886946E-2   9.145894E-2   -1.021446E-4   -8.855283E-6   8.855283E-6   -1.021446E-4   1.025277E-4   -1.750452E+2   -8.504521E+1   
5.278358E+3   5.000451E+1   5.000451E+1   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   -6.887407E-2   9.315256E-2   -1.032504E-4   -9.959111E-6   9.959111E-6   -1.032504E-4   1.037296E-4   -1.744905E+2   -8.449053E+1   
5.300541E+3   5.002068E+1   5.002068E+1   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   -7.023377E-2   9.191178E-2   -1.032830E-4   -8.142248E-6   8.142248E-6   -1.032830E-4   1.036034E-4   -1.754924E+2   -8.549245E+1   
5.322770E+3   5.001031E+1   5.001031E+1   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   -6.965208E-2   9.223300E-2   -1.031326E-4   -8.782490E-6   8.782490E-6   -1.031326E-4   1.035058E-4   -1.751326E+2   -8.513259E+1   
5.345047E+3   5.000240E+1   5.000240E+1   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   -6.871760E-2   9.290890E-2   -1.029950E-4   -9.915545E-6   9.915545E-6   -1.029950E-4   1.034712E-4   -1.745010E+2   -8.450096E+1   
5.367357E+3   5.000839E+1   5.000839E+1   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   -6.879124E-2   9.156234E-2   -1.021635E-4   -8.980737E-6   8.980737E-6   -1.021635E-4   1.025575E-4   -1.749763E+2   -8.497630E+1   
5.389576E+3   5.001040E+1   5.001040E+1   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   -6.859919E-2   9.313099E-2   -1.030665E-4   -1.014832E-5   1.014832E-5   -1.030665E-4   1.035649E-4   -1.743766E+2   -8.437656E+1   
5.411755E+3   5.002639E+1   5.002639E+1   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   -6.851820E-2   9.301354E-2   -1.029399E-4   -1.013144E-5   1.013144E-5   -1.029399E-4   1.034373E-4   -1.743790E+2   -8.437900E+1   
5.433826E+3   4.999581E+1   4.999581E+1   -7.000000E+0   -7.000000E+0   9.000000E+1   -6.000000E+0   -6.000000E+0   -6.912716E-2   9.318595E-2   -1.034287E-4   -9.793746E-6   9.793746E-6   -1.034287E-4   1.038913E-4   -1.745907E+2   -8.459074E+1   
5.454858E+3   5.003210E+1   5.003210E+1   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   -6.986929E-2   9.335532E-2   -1.039978E-4   -9.355579E-6   9.355579E-6   -1.039978E-4   1.044178E-4   -1.748595E+2   -8.485954E+1   
5.476934E+3   5.002691E+1   5.002691E+1   -3.000000E+0   -3.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   -6.948856E-2   9.330805E-2   -1.037316E-4   -9.606271E-6   9.606271E-6   -1.037316E-4   1.041755E-4   -1.747091E+2   -8.470910E+1   
5.497928E+3   5.003539E+1   5.003539E+1   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   -6.997606E-2   9.257266E-2   -1.035541E-4   -8.764923E-6   8.764923E-6   -1.035541E-4   1.039243E-4   -1.751620E+2   -8.516196E+1   
5.519913E+3   5.002349E+1   5.002349E+1   0.000000E+0   0.000000E+0   9.000000E+1   0.000000E+0   0.000000E+0   -7.036047E-2   9.276319E-2   -1.039158E-4   -8.605159E-6   8.605159E-6   -1.039158E-4   1.042715E-4   -1.752662E+2   -8.526620E+1   
5.541945E+3   5.000930E+1   5.000930E+1   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   -6.915171E-2   9.312428E-2   -1.034037E-4   -9.735272E-6   9.735272E-6   -1.034037E-4   1.038609E-4   -1.746216E+2   -8.462156E+1   
5.563418E+3   5.001599E+1   5.001599E+1   3.000000E+0   3.000000E+0   9.000000E+1   3.000000E+0   3.000000E+0   -7.078568E-2   9.226214E-2   -1.038524E-4   -7.963089E-6   7.963089E-6   -1.038524E-4   1.041572E-4   -1.756153E+2   -8.561531E+1   
5.585152E+3   5.003521E+1   5.003521E+1   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   -7.089153E-2   9.281897E-2   -1.042805E-4   -8.248844E-6   8.248844E-6   -1.042805E-4   1.046062E-4   -1.754772E+2   -8.547718E+1   
5.606672E+3   5.003939E+1   5.003939E+1   6.000000E+0   6.000000E+0   9.000000E+1   7.000000E+0   7.000000E+0   -7.010830E-2   9.227688E-2   -1.034432E-4   -8.473744E-6   8.473744E-6   -1.034432E-4   1.037897E-4   -1.753170E+2   -8.531696E+1   
5.628213E+3   5.002310E+1   5.002310E+1   9.000000E+0   9.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   -6.996257E-2   9.398182E-2   -1.044635E-4   -9.696169E-6   9.696169E-6   -1.044635E-4   1.049125E-4   -1.746971E+2   -8.469707E+1   
5.650195E+3   5.004061E+1   5.004061E+1   1.000000E+1   1.000000E+1   9.000000E+1   1.100000E+1   1.100000E+1   -6.899586E-2   9.268984E-2   -1.030244E-4   -9.566518E-6   9.566518E-6   -1.030244E-4   1.034676E-4   -1.746949E+2   -8.469491E+1   
5.672035E+3   4.999780E+1   4.999780E+1   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   -6.895812E-2   9.380447E-2   -1.037270E-4   -1.032315E-5   1.032315E-5   -1.037270E-4   1.042394E-4   -1.743165E+2   -8.431651E+1   
5.693900E+3   5.005361E+1   5.005361E+1   1.500000E+1   1.500000E+1   9.000000E+1   1.600000E+1   1.600000E+1   -7.018407E-2   9.305187E-2   -1.039948E-4   -8.924367E-6   8.924367E-6   -1.039948E-4   1.043770E-4   -1.750951E+2   -8.509515E+1   
5.715966E+3   5.001510E+1   5.001510E+1   1.600000E+1   1.600000E+1   9.000000E+1   1.800000E+1   1.800000E+1   -6.937353E-2   9.403335E-2   -1.041329E-4   -1.016553E-5   1.016553E-5   -1.041329E-4   1.046279E-4   -1.744244E+2   -8.442441E+1   
5.737910E+3   5.002529E+1   5.002529E+1   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   -7.070379E-2   9.338814E-2   -1.045351E-4   -8.759813E-6   8.759813E-6   -1.045351E-4   1.049015E-4   -1.752099E+2   -8.520993E+1   
5.759792E+3   4.999911E+1   4.999911E+1   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   -7.064243E-2   9.336971E-2   -1.044852E-4   -8.793139E-6   8.793139E-6   -1.044852E-4   1.048545E-4   -1.751895E+2   -8.518950E+1   
5.781658E+3   5.003079E+1   5.003079E+1   2.300000E+1   2.300000E+1   9.000000E+1   2.300000E+1   2.300000E+1   -6.953736E-2   9.320218E-2   -1.036928E-4   -9.500966E-6   9.500966E-6   -1.036928E-4   1.041272E-4   -1.747648E+2   -8.476483E+1   
5.803694E+3   5.000161E+1   5.000161E+1   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   -7.070623E-2   9.360354E-2   -1.046769E-4   -8.898830E-6   8.898830E-6   -1.046769E-4   1.050545E-4   -1.751408E+2   -8.514083E+1   
5.825600E+3   5.002300E+1   5.002300E+1   2.600000E+1   2.600000E+1   9.000000E+1   2.700000E+1   2.700000E+1   -7.078877E-2   9.386277E-2   -1.048968E-4   -9.007252E-6   9.007252E-6   -1.048968E-4   1.052828E-4   -1.750922E+2   -8.509218E+1   
5.847444E+3   5.003460E+1   5.003460E+1   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   -7.008590E-2   9.383486E-2   -1.044440E-4   -9.508870E-6   9.508870E-6   -1.044440E-4   1.048760E-4   -1.747980E+2   -8.479798E+1   
5.869345E+3   5.003109E+1   5.003109E+1   3.100000E+1   3.100000E+1   9.000000E+1   3.100000E+1   3.100000E+1   -7.085503E-2   9.374833E-2   -1.048632E-4   -8.883430E-6   8.883430E-6   -1.048632E-4   1.052388E-4   -1.751578E+2   -8.515778E+1   
5.891371E+3   5.000881E+1   5.000881E+1   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   -7.100567E-2   9.447886E-2   -1.054321E-4   -9.249608E-6   9.249608E-6   -1.054321E-4   1.058371E-4   -1.749863E+2   -8.498625E+1   
5.913312E+3   5.001489E+1   5.001489E+1   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   -7.112132E-2   9.481880E-2   -1.057250E-4   -9.386315E-6   9.386315E-6   -1.057250E-4   1.061408E-4   -1.749266E+2   -8.492656E+1   
5.935285E+3   5.001989E+1   5.001989E+1   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   -7.009387E-2   9.377226E-2   -1.044082E-4   -9.462049E-6   9.462049E-6   -1.044082E-4   1.048361E-4   -1.748217E+2   -8.482168E+1   
5.957242E+3   5.001611E+1   5.001611E+1   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   -7.119404E-2   9.470558E-2   -1.056962E-4   -9.258507E-6   9.258507E-6   -1.056962E-4   1.061010E-4   -1.749939E+2   -8.499393E+1   
5.979100E+3   5.002789E+1   5.002789E+1   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   -7.018101E-2   9.423554E-2   -1.047638E-4   -9.700479E-6   9.700479E-6   -1.047638E-4   1.052119E-4   -1.747098E+2   -8.470985E+1   
6.000958E+3   5.000839E+1   5.000839E+1   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   -7.080778E-2   9.500443E-2   -1.056521E-4   -9.739579E-6   9.739579E-6   -1.056521E-4   1.061000E-4   -1.747331E+2   -8.473305E+1   
6.022863E+3   5.000302E+1   5.000302E+1   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   -7.071021E-2   9.373882E-2   -1.047675E-4   -8.984322E-6   8.984322E-6   -1.047675E-4   1.051520E-4   -1.750986E+2   -8.509860E+1   
6.044834E+3   5.001370E+1   5.001370E+1   4.600000E+1   4.600000E+1   9.000000E+1   4.800000E+1   4.800000E+1   -7.010062E-2   9.449049E-2   -1.048801E-4   -9.926621E-6   9.926621E-6   -1.048801E-4   1.053489E-4   -1.745932E+2   -8.459322E+1   
6.066771E+3   5.003149E+1   5.003149E+1   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   -6.855162E-2   9.455954E-2   -1.039674E-4   -1.111745E-5   1.111745E-5   -1.039674E-4   1.045602E-4   -1.738964E+2   -8.389644E+1   
6.100681E+3   5.004131E+1   5.004131E+1   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   -7.249177E-2   9.580398E-2   -1.072139E-4   -9.016772E-6   9.016772E-6   -1.072139E-4   1.075924E-4   -1.751927E+2   -8.519269E+1   
6.123213E+3   5.003539E+1   5.003539E+1   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   -7.278261E-2   9.765369E-2   -1.085984E-4   -1.001094E-5   1.001094E-5   -1.085984E-4   1.090589E-4   -1.747332E+2   -8.473318E+1   
6.145537E+3   5.002770E+1   5.002770E+1   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   -7.475313E-2   9.882103E-2   -1.105770E-4   -9.316662E-6   9.316662E-6   -1.105770E-4   1.109688E-4   -1.751839E+2   -8.518392E+1   
6.167891E+3   5.003219E+1   5.003219E+1   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   -7.499889E-2   1.013754E-1   -1.123925E-4   -1.080488E-5   1.080488E-5   -1.123925E-4   1.129107E-4   -1.745087E+2   -8.450874E+1   
6.190487E+3   5.001760E+1   5.001760E+1   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   -7.458776E-2   1.016080E-1   -1.122898E-4   -1.126099E-5   1.126099E-5   -1.122898E-4   1.128531E-4   -1.742732E+2   -8.427324E+1   
6.212782E+3   5.001061E+1   5.001061E+1   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   -7.784990E-2   1.025032E-1   -1.148897E-4   -9.433470E-6   9.433470E-6   -1.148897E-4   1.152763E-4   -1.753060E+2   -8.530603E+1   
6.235169E+3   4.999740E+1   4.999740E+1   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   -7.834107E-2   1.037405E-1   -1.159992E-4   -9.879100E-6   9.879100E-6   -1.159992E-4   1.164191E-4   -1.751321E+2   -8.513214E+1   
6.257819E+3   5.002291E+1   5.002291E+1   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   -7.789806E-2   1.056496E-1   -1.169687E-4   -1.145493E-5   1.145493E-5   -1.169687E-4   1.175283E-4   -1.744068E+2   -8.440677E+1   
6.279912E+3   5.004470E+1   5.004470E+1   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   -8.031222E-2   1.070391E-1   -1.193662E-4   -1.057773E-5   1.057773E-5   -1.193662E-4   1.198340E-4   -1.749359E+2   -8.493592E+1   
6.302506E+3   5.000549E+1   5.000549E+1   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   -8.012445E-2   1.083178E-1   -1.200829E-4   -1.155260E-5   1.155260E-5   -1.200829E-4   1.206374E-4   -1.745048E+2   -8.450476E+1   
6.325862E+3   5.002401E+1   5.002401E+1   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   -8.072639E-2   1.096631E-1   -1.213312E-4   -1.198689E-5   1.198689E-5   -1.213312E-4   1.219219E-4   -1.743578E+2   -8.435779E+1   
6.348495E+3   5.000909E+1   5.000909E+1   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   -8.033306E-2   1.121527E-1   -1.227095E-4   -1.390546E-5   1.390546E-5   -1.227095E-4   1.234949E-4   -1.735348E+2   -8.353481E+1   
6.371145E+3   5.000680E+1   5.000680E+1   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   -8.346695E-2   1.128725E-1   -1.251158E-4   -1.205809E-5   1.205809E-5   -1.251158E-4   1.256955E-4   -1.744951E+2   -8.449510E+1   
6.394524E+3   5.001650E+1   5.001650E+1   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   -8.351327E-2   1.138622E-1   -1.257890E-4   -1.267086E-5   1.267086E-5   -1.257890E-4   1.264256E-4   -1.742479E+2   -8.424794E+1   
6.417118E+3   5.001730E+1   5.001730E+1   7.980000E+2   7.980000E+2   9.000000E+1   7.980000E+2   7.980000E+2   -8.500615E-2   1.150764E-1   -1.275028E-4   -1.236054E-5   1.236054E-5   -1.275028E-4   1.281006E-4   -1.744629E+2   -8.446286E+1   
6.439752E+3   4.999609E+1   4.999609E+1   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   -8.479352E-2   1.168500E-1   -1.285265E-4   -1.367733E-5   1.367733E-5   -1.285265E-4   1.292522E-4   -1.739257E+2   -8.392565E+1   
6.463010E+3   5.003271E+1   5.003271E+1   8.980000E+2   8.980000E+2   9.000000E+1   8.980000E+2   8.980000E+2   -8.463524E-2   1.178048E-1   -1.290505E-4   -1.441858E-5   1.441858E-5   -1.290505E-4   1.298534E-4   -1.736249E+2   -8.362488E+1   
6.485651E+3   5.003869E+1   5.003869E+1   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   -8.727703E-2   1.189644E-1   -1.314390E-4   -1.322279E-5   1.322279E-5   -1.314390E-4   1.321025E-4   -1.742554E+2   -8.425536E+1   
6.508289E+3   5.002270E+1   5.002270E+1   9.980000E+2   9.980000E+2   9.000000E+1   9.980000E+2   9.980000E+2   -8.812683E-2   1.219201E-1   -1.338894E-4   -1.452657E-5   1.452657E-5   -1.338894E-4   1.346751E-4   -1.738078E+2   -8.380781E+1   
6.531801E+3   5.002361E+1   5.002361E+1   1.048000E+3   1.048000E+3   9.000000E+1   1.048000E+3   1.048000E+3   -8.938808E-2   1.217452E-1   -1.345553E-4   -1.347938E-5   1.347938E-5   -1.345553E-4   1.352287E-4   -1.742793E+2   -8.427935E+1   
6.554621E+3   5.002340E+1   5.002340E+1   1.098000E+3   1.098000E+3   9.000000E+1   1.098000E+3   1.098000E+3   -8.938837E-2   1.232295E-1   -1.355221E-4   -1.444953E-5   1.444953E-5   -1.355221E-4   1.362903E-4   -1.739140E+2   -8.391405E+1   
6.577399E+3   5.000060E+1   5.000060E+1   1.148000E+3   1.148000E+3   9.000000E+1   1.148000E+3   1.148000E+3   -9.038207E-2   1.247429E-1   -1.371221E-4   -1.470399E-5   1.470399E-5   -1.371221E-4   1.379083E-4   -1.738794E+2   -8.387940E+1   
6.600670E+3   5.001711E+1   5.001711E+1   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   -9.132304E-2   1.263256E-1   -1.387347E-4   -1.504277E-5   1.504277E-5   -1.387347E-4   1.395479E-4   -1.738117E+2   -8.381169E+1   
6.623751E+3   5.001690E+1   5.001690E+1   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   -9.083063E-2   1.280483E-1   -1.395522E-4   -1.653319E-5   1.653319E-5   -1.395522E-4   1.405282E-4   -1.732435E+2   -8.324348E+1   
6.646287E+3   5.005432E+1   5.005432E+1   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   -9.358572E-2   1.288818E-1   -1.417984E-4   -1.504038E-5   1.504038E-5   -1.417984E-4   1.425939E-4   -1.739453E+2   -8.394535E+1   
6.669328E+3   5.001800E+1   5.001800E+1   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   -9.544956E-2   1.312113E-1   -1.444679E-4   -1.518478E-5   1.518478E-5   -1.444679E-4   1.452637E-4   -1.739998E+2   -8.399977E+1   
6.691866E+3   5.004391E+1   5.004391E+1   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   -9.476758E-2   1.324084E-1   -1.448259E-4   -1.647182E-5   1.647182E-5   -1.448259E-4   1.457596E-4   -1.735113E+2   -8.351133E+1   
6.714391E+3   5.003329E+1   5.003329E+1   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   -9.662036E-2   1.343525E-1   -1.472376E-4   -1.637248E-5   1.637248E-5   -1.472376E-4   1.481451E-4   -1.736549E+2   -8.365491E+1   
6.737178E+3   5.001351E+1   5.001351E+1   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   -9.631691E-2   1.345403E-1   -1.471723E-4   -1.671967E-5   1.671967E-5   -1.471723E-4   1.481190E-4   -1.735186E+2   -8.351864E+1   
6.759727E+3   5.000839E+1   5.000839E+1   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   -9.879315E-2   1.368658E-1   -1.502178E-4   -1.640850E-5   1.640850E-5   -1.502178E-4   1.511113E-4   -1.737662E+2   -8.376622E+1   
6.782316E+3   4.999639E+1   4.999639E+1   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   -9.816299E-2   1.376484E-1   -1.503379E-4   -1.738625E-5   1.738625E-5   -1.503379E-4   1.513399E-4   -1.734032E+2   -8.340317E+1   
6.805375E+3   5.003060E+1   5.003060E+1   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   -9.971534E-2   1.397570E-1   -1.526709E-4   -1.761661E-5   1.761661E-5   -1.526709E-4   1.536840E-4   -1.734178E+2   -8.341778E+1   
6.827971E+3   5.002331E+1   5.002331E+1   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   -1.003372E-1   1.413106E-1   -1.540673E-4   -1.817236E-5   1.817236E-5   -1.540673E-4   1.551353E-4   -1.732730E+2   -8.327300E+1   
6.850786E+3   5.003201E+1   5.003201E+1   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   -1.020583E-1   1.416091E-1   -1.553257E-4   -1.709453E-5   1.709453E-5   -1.553257E-4   1.562636E-4   -1.737195E+2   -8.371953E+1   
6.873584E+3   5.000729E+1   5.000729E+1   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   -1.020090E-1   1.435732E-1   -1.565744E-4   -1.841511E-5   1.841511E-5   -1.565744E-4   1.576536E-4   -1.732921E+2   -8.329211E+1   
6.896168E+3   4.998541E+1   4.998541E+1   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   -1.018644E-1   1.447838E-1   -1.572735E-4   -1.931346E-5   1.931346E-5   -1.572735E-4   1.584549E-4   -1.729990E+2   -8.299903E+1   
6.918711E+3   5.003521E+1   5.003521E+1   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   -1.028879E-1   1.461168E-1   -1.587745E-4   -1.942795E-5   1.942795E-5   -1.587745E-4   1.599587E-4   -1.730239E+2   -8.302386E+1   
6.941502E+3   5.002850E+1   5.002850E+1   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   -1.052266E-1   1.478183E-1   -1.613285E-4   -1.881057E-5   1.881057E-5   -1.613285E-4   1.624214E-4   -1.733495E+2   -8.334946E+1   
6.964038E+3   5.001159E+1   5.001159E+1   1.999000E+3   1.999000E+3   9.000000E+1   2.000000E+3   2.000000E+3   -1.054380E-1   1.499615E-1   -1.628550E-4   -2.005543E-5   2.005543E-5   -1.628550E-4   1.640853E-4   -1.729794E+2   -8.297943E+1   
7.002016E+3   5.002520E+1   5.002520E+1   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   -1.143181E-1   1.638798E-1   -1.774099E-4   -2.258678E-5   2.258678E-5   -1.774099E-4   1.788420E-4   -1.727445E+2   -8.274447E+1   
7.028660E+3   5.000759E+1   5.000759E+1   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   -1.261744E-1   1.812464E-1   -1.960508E-4   -2.517129E-5   2.517129E-5   -1.960508E-4   1.976600E-4   -1.726837E+2   -8.268372E+1   
7.054613E+3   5.001559E+1   5.001559E+1   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -1.351045E-1   1.950982E-1   -2.105933E-4   -2.762221E-5   2.762221E-5   -2.105933E-4   2.123971E-4   -1.725275E+2   -8.252753E+1   
7.080410E+3   5.001251E+1   5.001251E+1   3.999000E+3   3.999000E+3   9.000000E+1   4.000000E+3   4.000000E+3   -1.449022E-1   2.123893E-1   -2.279123E-4   -3.167995E-5   3.167995E-5   -2.279123E-4   2.301035E-4   -1.720866E+2   -8.208656E+1   
7.106861E+3   5.001541E+1   5.001541E+1   4.498000E+3   4.498000E+3   9.000000E+1   4.499000E+3   4.499000E+3   -1.542026E-1   2.251632E-1   -2.419817E-4   -3.315232E-5   3.315232E-5   -2.419817E-4   2.442421E-4   -1.721988E+2   -8.219885E+1   
7.132804E+3   5.002542E+1   5.002542E+1   4.997000E+3   4.997000E+3   9.000000E+1   4.999000E+3   4.999000E+3   -1.586484E-1   2.354432E-1   -2.514255E-4   -3.658489E-5   3.658489E-5   -2.514255E-4   2.540733E-4   -1.717210E+2   -8.172100E+1   
7.158417E+3   5.000161E+1   5.000161E+1   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -1.610260E-1   2.403154E-1   -2.560687E-4   -3.801159E-5   3.801159E-5   -2.560687E-4   2.588746E-4   -1.715565E+2   -8.155650E+1   
7.184910E+3   5.000759E+1   5.000759E+1   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -1.490243E-1   2.291709E-1   -2.413903E-4   -3.960244E-5   3.960244E-5   -2.413903E-4   2.446173E-4   -1.706831E+2   -8.068307E+1   
7.210810E+3   4.999230E+1   4.999230E+1   6.498000E+3   6.498000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -1.298740E-1   2.118310E-1   -2.182574E-4   -4.243028E-5   4.243028E-5   -2.182574E-4   2.223435E-4   -1.689987E+2   -7.899865E+1   
7.236960E+3   5.002831E+1   5.002831E+1   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -1.145095E-1   1.958369E-1   -1.983416E-4   -4.333784E-5   4.333784E-5   -1.983416E-4   2.030211E-4   -1.676745E+2   -7.767453E+1   
7.262619E+3   5.002459E+1   5.002459E+1   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -1.008409E-1   1.810780E-1   -1.802787E-4   -4.379856E-5   4.379856E-5   -1.802787E-4   1.855229E-4   -1.663446E+2   -7.634460E+1   
7.288063E+3   5.004781E+1   5.004781E+1   7.999000E+3   7.999000E+3   9.000000E+1   8.000000E+3   8.000000E+3   -9.398181E-2   1.771980E-1   -1.735111E-4   -4.633516E-5   4.633516E-5   -1.735111E-4   1.795913E-4   -1.650484E+2   -7.504838E+1   
7.314512E+3   4.999371E+1   4.999371E+1   8.498000E+3   8.498000E+3   9.000000E+1   8.499000E+3   8.499000E+3   -8.931479E-2   1.762527E-1   -1.700101E-4   -4.916907E-5   4.916907E-5   -1.700101E-4   1.769775E-4   -1.638695E+2   -7.386946E+1   
7.340951E+3   5.004391E+1   5.004391E+1   8.998000E+3   8.998000E+3   9.000000E+1   8.999000E+3   8.999000E+3   -9.227235E-2   1.826843E-1   -1.760275E-4   -5.118638E-5   5.118638E-5   -1.760275E-4   1.833186E-4   -1.637863E+2   -7.378629E+1   
7.367334E+3   5.000030E+1   5.000030E+1   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -9.859427E-2   1.940118E-1   -1.873134E-4   -5.391604E-5   5.391604E-5   -1.873134E-4   1.949186E-4   -1.639421E+2   -7.394214E+1   
7.393235E+3   5.001141E+1   5.001141E+1   9.999000E+3   9.999000E+3   9.000000E+1   1.000000E+4   1.000000E+4   -1.081208E-1   2.089186E-1   -2.029118E-4   -5.661554E-5   5.661554E-5   -2.029118E-4   2.106621E-4   -1.644101E+2   -7.441007E+1   
@@END Data.
@Time at end of measurement: 15:16:01
@NO Instrument  Changes.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -9499.000      -9999.000      250.000        Coercive Field: Field at which M//H changes sign
Ms  emu                                 3.047E-4       -2.561E-4      2.804E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -1.039E-4      1.421E-4       1.230E-4       Remanent Magnetization: M at H=0        
S                                       0.341          0.555          0.448          Squareness: Mr/Ms                       
S*                                      1.427          1.317          1.372          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
