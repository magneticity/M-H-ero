@Filename: c:\vsm-lv\Will\data\AJA335e-FePtFeRh_1030nm_Tann_6\AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_120deg.VHD
@Measurement Controlfilename: C:\vsm-lv\Will\Recipes\10kOe OoP loop 120deg.VHC
@Signal Manipulation filename: c:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA335e-FePtFeRh_1030nm_Tann_6
@Date: 08 November 2019    (2019-08-11)
@Time: 13:09:33
@Test ID: AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_120deg
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 90.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Sample Temperature to 120.0106 [degC] and wait 60.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Applied Field to 9999.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 3:      Set Auto Range Signal to 12.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 5
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 5.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 10000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To: 50.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: 50.0000 [Oe] To: -50.0000 [Oe] Min Stepsize/Sweeprate =  2.0000 [Oe] Max Stepsize/Sweeprate =  2.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -50.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -10000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 4 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 20 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.706
@Y Coils Correction Factor: 0.964
@Sample Shape Correction Factor: 0.919
@Coil Angle Alpha: 42.300
@Coil Angle Beta: -47.320
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
15000.000000   1.000000
15249.000000   1.000524
15499.000000   1.000702
15750.000000   1.001233
16000.000000   1.001406
16250.000000   1.001585
16499.000000   1.001758
16749.000000   1.001937
16999.000000   1.002110
17249.000000   1.001937
17499.000000   1.002289
17749.000000   1.002289
17999.000000   1.002289
18249.000000   1.002462
18499.000000   1.002462
18748.000000   1.002462
18999.000000   1.002462
19249.000000   1.002462
19499.000000   1.002642
19749.000000   1.002642
19999.000000   1.002462
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = No
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 25 October 2019  12:02:56
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 5
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 13:09:33
@@Data
New Section: Section 0: 
2.967200E+1   1.200115E+2   1.200115E+2   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -2.015586E-1   2.867262E-1   -3.113547E-4   -3.837447E-5   3.837447E-5   -3.113547E-4   3.137106E-4   -1.729737E+2   -8.297373E+1   
5.506100E+1   1.200159E+2   1.200159E+2   9.498000E+3   9.498000E+3   9.000000E+1   9.498000E+3   9.498000E+3   -1.827857E-1   2.660381E-1   -2.862745E-4   -3.873417E-5   3.873417E-5   -2.862745E-4   2.888830E-4   -1.722944E+2   -8.229443E+1   
8.016800E+1   1.200712E+2   1.200712E+2   8.997000E+3   8.997000E+3   9.000000E+1   8.998000E+3   8.998000E+3   -1.654089E-1   2.421811E-1   -2.599935E-4   -3.598960E-5   3.598960E-5   -2.599935E-4   2.624726E-4   -1.721189E+2   -8.211891E+1   
1.055250E+2   1.200067E+2   1.200067E+2   8.498000E+3   8.498000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -1.536219E-1   2.260174E-1   -2.421789E-4   -3.414025E-5   3.414025E-5   -2.421789E-4   2.445735E-4   -1.719758E+2   -8.197582E+1   
1.309210E+2   1.200252E+2   1.200252E+2   7.998000E+3   7.998000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -1.351413E-1   2.014562E-1   -2.147569E-4   -3.175165E-5   3.175165E-5   -2.147569E-4   2.170915E-4   -1.715898E+2   -8.158979E+1   
1.565640E+2   1.200996E+2   1.200996E+2   7.498000E+3   7.498000E+3   9.000000E+1   7.498000E+3   7.498000E+3   -1.202993E-1   1.810305E-1   -1.922779E-4   -2.937551E-5   2.937551E-5   -1.922779E-4   1.945089E-4   -1.713137E+2   -8.131373E+1   
1.815120E+2   1.200591E+2   1.200591E+2   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -1.047213E-1   1.587607E-1   -1.681427E-4   -2.633812E-5   2.633812E-5   -1.681427E-4   1.701930E-4   -1.710974E+2   -8.109745E+1   
2.068970E+2   1.199903E+2   1.199903E+2   6.497000E+3   6.497000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -8.997375E-2   1.395726E-1   -1.465282E-4   -2.470126E-5   2.470126E-5   -1.465282E-4   1.485956E-4   -1.704312E+2   -8.043122E+1   
2.319970E+2   1.200180E+2   1.200180E+2   5.998000E+3   5.998000E+3   9.000000E+1   5.998000E+3   5.998000E+3   -7.707554E-2   1.196612E-1   -1.255858E-4   -2.122363E-5   2.122363E-5   -1.255858E-4   1.273665E-4   -1.704078E+2   -8.040781E+1   
2.578540E+2   1.200206E+2   1.200206E+2   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -6.014336E-2   9.866731E-2   -1.014444E-4   -2.002200E-5   2.002200E-5   -1.014444E-4   1.034014E-4   -1.688351E+2   -7.883508E+1   
2.831530E+2   1.199954E+2   1.199954E+2   4.997000E+3   4.997000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -4.560065E-2   7.874143E-2   -7.947591E-5   -1.775126E-5   1.775126E-5   -7.947591E-5   8.143420E-5   -1.674094E+2   -7.740941E+1   
3.082950E+2   1.200413E+2   1.200413E+2   4.498000E+3   4.498000E+3   9.000000E+1   4.498000E+3   4.498000E+3   -3.183849E-2   5.941749E-2   -5.838202E-5   -1.529674E-5   1.529674E-5   -5.838202E-5   6.035272E-5   -1.653179E+2   -7.531790E+1   
3.345640E+2   1.200141E+2   1.200141E+2   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -1.768454E-2   3.975775E-2   -3.682721E-5   -1.291246E-5   1.291246E-5   -3.682721E-5   3.902531E-5   -1.606782E+2   -7.067817E+1   
3.599700E+2   1.200954E+2   1.200954E+2   3.498000E+3   3.498000E+3   9.000000E+1   3.498000E+3   3.498000E+3   -2.545778E-3   2.030149E-2   -1.479606E-5   -1.138960E-5   1.138960E-5   -1.479606E-5   1.867208E-5   -1.424119E+2   -5.241191E+1   
3.852760E+2   1.200839E+2   1.200839E+2   2.998000E+3   2.998000E+3   9.000000E+1   2.998000E+3   2.998000E+3   1.088813E-2   1.525074E-3   5.738289E-6   -9.050252E-6   9.050252E-6   5.738289E-6   1.071611E-5   -5.762337E+1   3.237663E+1   
4.109630E+2   1.199443E+2   1.199443E+2   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   2.664695E-2   -1.944552E-2   2.913905E-5   -6.995976E-6   6.995976E-6   2.913905E-5   2.996712E-5   -1.350057E+1   7.649943E+1   
4.367610E+2   1.200055E+2   1.200055E+2   1.999000E+3   1.999000E+3   9.000000E+1   1.999000E+3   1.999000E+3   4.182981E-2   -4.059499E-2   5.230023E-5   -4.398769E-6   4.398769E-6   5.230023E-5   5.248489E-5   -4.807610E+0   8.519239E+1   
4.706080E+2   1.200428E+2   1.200428E+2   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   4.360769E-2   -4.202524E-2   5.433091E-5   -4.778687E-6   4.778687E-6   5.433091E-5   5.454066E-5   -5.026527E+0   8.497347E+1   
4.929300E+2   1.200708E+2   1.200708E+2   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   4.440444E-2   -4.262994E-2   5.521733E-5   -4.972654E-6   4.972654E-6   5.521733E-5   5.544078E-5   -5.145949E+0   8.485405E+1   
5.152260E+2   1.200564E+2   1.200564E+2   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   4.554112E-2   -4.480513E-2   5.733675E-5   -4.391297E-6   4.391297E-6   5.733675E-5   5.750467E-5   -4.379609E+0   8.562039E+1   
5.374520E+2   1.200157E+2   1.200157E+2   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   4.684011E-2   -4.701776E-2   5.958092E-5   -3.905515E-6   3.905515E-6   5.958092E-5   5.970878E-5   -3.750359E+0   8.624964E+1   
5.597190E+2   1.200398E+2   1.200398E+2   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   4.997255E-2   -4.822473E-2   6.230362E-5   -5.433279E-6   5.433279E-6   6.230362E-5   6.254008E-5   -4.983954E+0   8.501605E+1   
5.819800E+2   1.200796E+2   1.200796E+2   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   5.078216E-2   -5.087329E-2   6.452914E-5   -4.300546E-6   4.300546E-6   6.452914E-5   6.467229E-5   -3.812840E+0   8.618716E+1   
6.045170E+2   1.200455E+2   1.200455E+2   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   5.257723E-2   -5.352922E-2   6.736871E-5   -3.891861E-6   3.891861E-6   6.736871E-5   6.748104E-5   -3.306277E+0   8.669372E+1   
6.267680E+2   1.199999E+2   1.199999E+2   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   5.426061E-2   -5.536998E-2   6.960833E-5   -3.933503E-6   3.933503E-6   6.960833E-5   6.971938E-5   -3.234293E+0   8.676571E+1   
6.488110E+2   1.200238E+2   1.200238E+2   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   5.560437E-2   -5.732425E-2   7.171190E-5   -3.649744E-6   3.649744E-6   7.171190E-5   7.180472E-5   -2.913528E+0   8.708647E+1   
6.710290E+2   1.199886E+2   1.199886E+2   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   5.637870E-2   -5.946413E-2   7.358430E-5   -2.823468E-6   2.823468E-6   7.358430E-5   7.363845E-5   -2.197391E+0   8.780261E+1   
6.933170E+2   1.200577E+2   1.200577E+2   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   5.891128E-2   -6.029185E-2   7.568915E-5   -4.155498E-6   4.155498E-6   7.568915E-5   7.580314E-5   -3.142507E+0   8.685749E+1   
7.156150E+2   1.199942E+2   1.199942E+2   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   5.951106E-2   -6.325457E-2   7.798955E-5   -2.662182E-6   2.662182E-6   7.798955E-5   7.803497E-5   -1.955039E+0   8.804496E+1   
7.378890E+2   1.199602E+2   1.199602E+2   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   6.090082E-2   -6.634580E-2   8.086205E-5   -1.669133E-6   1.669133E-6   8.086205E-5   8.087928E-5   -1.182517E+0   8.881748E+1   
7.601990E+2   1.200357E+2   1.200357E+2   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   6.104993E-2   -6.712934E-2   8.146455E-5   -1.267155E-6   1.267155E-6   8.146455E-5   8.147441E-5   -8.911457E-1   8.910885E+1   
7.824820E+2   1.199828E+2   1.199828E+2   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   6.387181E-2   -6.829148E-2   8.396606E-5   -2.594533E-6   2.594533E-6   8.396606E-5   8.400613E-5   -1.769864E+0   8.823014E+1   
8.047290E+2   1.200521E+2   1.200521E+2   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   6.513210E-2   -7.102652E-2   8.652653E-5   -1.738593E-6   1.738593E-6   8.652653E-5   8.654400E-5   -1.151100E+0   8.884890E+1   
8.269910E+2   1.200404E+2   1.200404E+2   1.148000E+3   1.148000E+3   9.000000E+1   1.148000E+3   1.148000E+3   6.775672E-2   -7.319709E-2   8.956286E-5   -2.260789E-6   2.260789E-6   8.956286E-5   8.959139E-5   -1.445981E+0   8.855402E+1   
8.493050E+2   1.199625E+2   1.199625E+2   1.097000E+3   1.097000E+3   9.000000E+1   1.098000E+3   1.098000E+3   6.732599E-2   -7.541243E-2   9.073939E-5   -4.938717E-7   4.938717E-7   9.073939E-5   9.074074E-5   -3.118434E-1   8.968816E+1   
8.716340E+2   1.200142E+2   1.200142E+2   1.047000E+3   1.047000E+3   9.000000E+1   1.048000E+3   1.048000E+3   6.884275E-2   -7.721176E-2   9.284901E-5   -4.393684E-7   4.393684E-7   9.284901E-5   9.285005E-5   -2.711258E-1   8.972887E+1   
8.938050E+2   1.199911E+2   1.199911E+2   9.980000E+2   9.980000E+2   9.000000E+1   9.980000E+2   9.980000E+2   6.930601E-2   -7.924120E-2   9.445717E-5   5.447776E-7   -5.447776E-7   9.445717E-5   9.445874E-5   3.304473E-1   9.033045E+1   
9.156420E+2   1.200303E+2   1.200303E+2   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   7.116886E-2   -8.047081E-2   9.640970E-5   -2.915480E-8   2.915480E-8   9.640970E-5   9.640971E-5   -1.732654E-2   8.998267E+1   
9.374790E+2   1.200271E+2   1.200271E+2   8.970000E+2   8.970000E+2   9.000000E+1   8.980000E+2   8.980000E+2   7.326211E-2   -8.056593E-2   9.776580E-5   -1.515200E-6   1.515200E-6   9.776580E-5   9.777754E-5   -8.879138E-1   8.911209E+1   
9.593560E+2   1.200456E+2   1.200456E+2   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   7.423864E-2   -8.414466E-2   1.007003E-4   1.021997E-7   -1.021997E-7   1.007003E-4   1.007004E-4   5.814886E-2   9.005815E+1   
9.811850E+2   1.200230E+2   1.200230E+2   7.980000E+2   7.980000E+2   9.000000E+1   7.980000E+2   7.980000E+2   7.591125E-2   -8.567279E-2   1.027297E-4   -1.358652E-7   1.358652E-7   1.027297E-4   1.027298E-4   -7.577651E-2   8.992422E+1   
1.003084E+3   1.199516E+2   1.199516E+2   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   7.702954E-2   -8.750465E-2   1.046141E-4   2.346271E-7   -2.346271E-7   1.046141E-4   1.046144E-4   1.285020E-1   9.012850E+1   
1.024957E+3   1.200302E+2   1.200302E+2   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   7.782504E-2   -8.922668E-2   1.062275E-4   7.720664E-7   -7.720664E-7   1.062275E-4   1.062303E-4   4.164212E-1   9.041642E+1   
1.046828E+3   1.200113E+2   1.200113E+2   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   7.913444E-2   -9.006669E-2   1.075841E-4   3.527629E-7   -3.527629E-7   1.075841E-4   1.075847E-4   1.878693E-1   9.018787E+1   
1.068658E+3   1.200238E+2   1.200238E+2   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   8.017383E-2   -9.352958E-2   1.104820E-4   1.847943E-6   -1.847943E-6   1.104820E-4   1.104975E-4   9.582503E-1   9.095825E+1   
1.090554E+3   1.200465E+2   1.200465E+2   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   8.166394E-2   -9.502404E-2   1.123766E-4   1.722843E-6   -1.722843E-6   1.123766E-4   1.123898E-4   8.783312E-1   9.087833E+1   
1.112380E+3   1.199301E+2   1.199301E+2   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   8.305064E-2   -9.679773E-2   1.143891E-4   1.856786E-6   -1.856786E-6   1.143891E-4   1.144042E-4   9.299543E-1   9.092995E+1   
1.134463E+3   1.199704E+2   1.199704E+2   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   8.511259E-2   -9.723644E-2   1.159496E-4   6.185241E-7   -6.185241E-7   1.159496E-4   1.159513E-4   3.056369E-1   9.030564E+1   
1.156340E+3   1.201286E+2   1.201286E+2   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   8.583049E-2   -1.002418E-1   1.183509E-4   2.052376E-6   -2.052376E-6   1.183509E-4   1.183687E-4   9.934926E-1   9.099349E+1   
1.178171E+3   1.199561E+2   1.199561E+2   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   8.650420E-2   -1.010266E-1   1.192785E-4   2.067133E-6   -2.067133E-6   1.192785E-4   1.192964E-4   9.928541E-1   9.099285E+1   
1.199995E+3   1.200724E+2   1.200724E+2   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   8.741139E-2   -1.039439E-1   1.217394E-4   3.303408E-6   -3.303408E-6   1.217394E-4   1.217842E-4   1.554345E+0   9.155434E+1   
1.222076E+3   1.200073E+2   1.200073E+2   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   8.981450E-2   -1.058494E-1   1.244661E-4   2.771734E-6   -2.771734E-6   1.244661E-4   1.244970E-4   1.275708E+0   9.127571E+1   
1.243860E+3   1.200445E+2   1.200445E+2   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   9.030662E-2   -1.071446E-1   1.256139E-4   3.254557E-6   -3.254557E-6   1.256139E-4   1.256561E-4   1.484156E+0   9.148416E+1   
1.265691E+3   1.199463E+2   1.199463E+2   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   9.169950E-2   -1.080074E-1   1.270370E-4   2.788361E-6   -2.788361E-6   1.270370E-4   1.270676E-4   1.257395E+0   9.125740E+1   
1.287468E+3   1.200076E+2   1.200076E+2   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   9.399502E-2   -1.105099E-1   1.300860E-4   2.726584E-6   -2.726584E-6   1.300860E-4   1.301146E-4   1.200735E+0   9.120074E+1   
1.309202E+3   1.200185E+2   1.200185E+2   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   9.620370E-2   -1.119033E-1   1.323591E-4   2.003979E-6   -2.003979E-6   1.323591E-4   1.323742E-4   8.674188E-1   9.086742E+1   
1.342343E+3   1.200082E+2   1.200082E+2   4.700000E+1   4.700000E+1   9.000000E+1   4.700000E+1   4.700000E+1   9.424935E-2   -1.125003E-1   1.315396E-4   3.839783E-6   -3.839783E-6   1.315396E-4   1.315956E-4   1.672051E+0   9.167205E+1   
1.363771E+3   1.200817E+2   1.200817E+2   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   9.579413E-2   -1.131467E-1   1.329157E-4   3.119824E-6   -3.119824E-6   1.329157E-4   1.329523E-4   1.344612E+0   9.134461E+1   
1.382860E+3   1.199918E+2   1.199918E+2   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   9.432176E-2   -1.129295E-1   1.318639E-4   4.066829E-6   -4.066829E-6   1.318639E-4   1.319266E-4   1.766505E+0   9.176651E+1   
1.405314E+3   1.200129E+2   1.200129E+2   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   9.457240E-2   -1.136520E-1   1.324894E-4   4.353802E-6   -4.353802E-6   1.324894E-4   1.325610E-4   1.882148E+0   9.188215E+1   
1.424372E+3   1.200094E+2   1.200094E+2   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   9.575610E-2   -1.131710E-1   1.329080E-4   3.163806E-6   -3.163806E-6   1.329080E-4   1.329456E-4   1.363639E+0   9.136364E+1   
1.446780E+3   1.200167E+2   1.200167E+2   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   9.589634E-2   -1.121046E-1   1.323001E-4   2.362892E-6   -2.362892E-6   1.323001E-4   1.323212E-4   1.023199E+0   9.102320E+1   
1.465882E+3   1.199931E+2   1.199931E+2   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   9.536246E-2   -1.128771E-1   1.324732E-4   3.262804E-6   -3.262804E-6   1.324732E-4   1.325134E-4   1.410905E+0   9.141091E+1   
1.488270E+3   1.201078E+2   1.201078E+2   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   9.617365E-2   -1.128443E-1   1.329533E-4   2.641369E-6   -2.641369E-6   1.329533E-4   1.329795E-4   1.138139E+0   9.113814E+1   
1.507306E+3   1.200271E+2   1.200271E+2   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   9.592668E-2   -1.123972E-1   1.325095E-4   2.531788E-6   -2.531788E-6   1.325095E-4   1.325337E-4   1.094587E+0   9.109459E+1   
1.529694E+3   1.200009E+2   1.200009E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   9.542169E-2   -1.131749E-1   1.327038E-4   3.413741E-6   -3.413741E-6   1.327038E-4   1.327477E-4   1.473581E+0   9.147358E+1   
1.548772E+3   1.199194E+2   1.199194E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   9.544225E-2   -1.130351E-1   1.326254E-4   3.307077E-6   -3.307077E-6   1.326254E-4   1.326666E-4   1.428401E+0   9.142840E+1   
1.571158E+3   1.200411E+2   1.200411E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   9.469764E-2   -1.132323E-1   1.322935E-4   3.986781E-6   -3.986781E-6   1.322935E-4   1.323536E-4   1.726136E+0   9.172614E+1   
1.590177E+3   1.200875E+2   1.200875E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   9.456720E-2   -1.127804E-1   1.319186E-4   3.787816E-6   -3.787816E-6   1.319186E-4   1.319729E-4   1.644698E+0   9.164470E+1   
1.612623E+3   1.200562E+2   1.200562E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   9.553240E-2   -1.141868E-1   1.334312E-4   3.993348E-6   -3.993348E-6   1.334312E-4   1.334910E-4   1.714244E+0   9.171424E+1   
1.631701E+3   1.200270E+2   1.200270E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   9.700600E-2   -1.134324E-1   1.338509E-4   2.410229E-6   -2.410229E-6   1.338509E-4   1.338726E-4   1.031603E+0   9.103160E+1   
1.654084E+3   1.199852E+2   1.199852E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.800000E+1   1.800000E+1   9.606320E-2   -1.136747E-1   1.334259E-4   3.265995E-6   -3.265995E-6   1.334259E-4   1.334659E-4   1.402204E+0   9.140220E+1   
1.673140E+3   1.200480E+2   1.200480E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   9.518264E-2   -1.134606E-1   1.327420E-4   3.777289E-6   -3.777289E-6   1.327420E-4   1.327958E-4   1.629961E+0   9.162996E+1   
1.695533E+3   1.200371E+2   1.200371E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   9.577726E-2   -1.131765E-1   1.329246E-4   3.151759E-6   -3.151759E-6   1.329246E-4   1.329620E-4   1.358279E+0   9.135828E+1   
1.714625E+3   1.200498E+2   1.200498E+2   1.300000E+1   1.300000E+1   9.000000E+1   1.300000E+1   1.300000E+1   9.584385E-2   -1.141239E-1   1.335828E-4   3.721875E-6   -3.721875E-6   1.335828E-4   1.336347E-4   1.595958E+0   9.159596E+1   
1.736394E+3   1.200831E+2   1.200831E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   9.543213E-2   -1.146497E-1   1.336708E-4   4.370173E-6   -4.370173E-6   1.336708E-4   1.337422E-4   1.872536E+0   9.187254E+1   
1.755066E+3   1.199851E+2   1.199851E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   9.595952E-2   -1.134345E-1   1.332053E-4   3.185622E-6   -3.185622E-6   1.332053E-4   1.332434E-4   1.369974E+0   9.136997E+1   
1.777095E+3   1.200895E+2   1.200895E+2   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   9.708883E-2   -1.140803E-1   1.343242E-4   2.772568E-6   -2.772568E-6   1.343242E-4   1.343528E-4   1.182467E+0   9.118247E+1   
1.795772E+3   1.199683E+2   1.199683E+2   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   9.624300E-2   -1.157959E-1   1.349186E-4   4.519777E-6   -4.519777E-6   1.349186E-4   1.349943E-4   1.918693E+0   9.191869E+1   
1.817778E+3   1.200274E+2   1.200274E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   9.584875E-2   -1.149019E-1   1.340926E-4   4.226905E-6   -4.226905E-6   1.340926E-4   1.341592E-4   1.805496E+0   9.180550E+1   
1.836496E+3   1.199920E+2   1.199920E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   9.564624E-2   -1.146454E-1   1.338003E-4   4.209003E-6   -4.209003E-6   1.338003E-4   1.338665E-4   1.801779E+0   9.180178E+1   
1.858526E+3   1.200872E+2   1.200872E+2   -1.000000E+0   -1.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   9.726679E-2   -1.150933E-1   1.350939E-4   3.303232E-6   -3.303232E-6   1.350939E-4   1.351343E-4   1.400681E+0   9.140068E+1   
1.880226E+3   1.199983E+2   1.199983E+2   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   9.629698E-2   -1.151713E-1   1.345451E-4   4.071484E-6   -4.071484E-6   1.345451E-4   1.346067E-4   1.733305E+0   9.173330E+1   
1.902268E+3   1.200388E+2   1.200388E+2   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   9.628259E-2   -1.162239E-1   1.352218E-4   4.770286E-6   -4.770286E-6   1.352218E-4   1.353059E-4   2.020414E+0   9.202041E+1   
1.924304E+3   1.200717E+2   1.200717E+2   -8.000000E+0   -8.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   9.768833E-2   -1.149556E-1   1.352648E-4   2.901378E-6   -2.901378E-6   1.352648E-4   1.352960E-4   1.228784E+0   9.122878E+1   
1.946388E+3   1.200932E+2   1.200932E+2   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   9.647367E-2   -1.148092E-1   1.344186E-4   3.704118E-6   -3.704118E-6   1.344186E-4   1.344696E-4   1.578477E+0   9.157848E+1   
1.968584E+3   1.200439E+2   1.200439E+2   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   9.787395E-2   -1.152789E-1   1.355902E-4   2.975499E-6   -2.975499E-6   1.355902E-4   1.356228E-4   1.257142E+0   9.125714E+1   
1.990784E+3   1.200561E+2   1.200561E+2   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   9.722230E-2   -1.153685E-1   1.352457E-4   3.516046E-6   -3.516046E-6   1.352457E-4   1.352914E-4   1.489210E+0   9.148921E+1   
2.013055E+3   1.200410E+2   1.200410E+2   -1.500000E+1   -1.500000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   9.729716E-2   -1.150611E-1   1.350918E-4   3.259713E-6   -3.259713E-6   1.350918E-4   1.351311E-4   1.382258E+0   9.138226E+1   
2.034983E+3   1.200104E+2   1.200104E+2   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   9.762698E-2   -1.159431E-1   1.358701E-4   3.592411E-6   -3.592411E-6   1.358701E-4   1.359176E-4   1.514550E+0   9.151455E+1   
2.057270E+3   1.199939E+2   1.199939E+2   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   9.724442E-2   -1.154066E-1   1.352841E-4   3.524562E-6   -3.524562E-6   1.352841E-4   1.353300E-4   1.492391E+0   9.149239E+1   
2.079514E+3   1.200397E+2   1.200397E+2   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   9.800988E-2   -1.161732E-1   1.362567E-4   3.459628E-6   -3.459628E-6   1.362567E-4   1.363006E-4   1.454457E+0   9.145446E+1   
2.101791E+3   1.200046E+2   1.200046E+2   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   9.803625E-2   -1.159247E-1   1.361112E-4   3.277663E-6   -3.277663E-6   1.361112E-4   1.361506E-4   1.379460E+0   9.137946E+1   
2.124066E+3   1.200671E+2   1.200671E+2   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   9.731775E-2   -1.157784E-1   1.355716E-4   3.713410E-6   -3.713410E-6   1.355716E-4   1.356225E-4   1.568983E+0   9.156898E+1   
2.146357E+3   1.200241E+2   1.200241E+2   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   9.834549E-2   -1.167037E-1   1.368097E-4   3.558198E-6   -3.558198E-6   1.368097E-4   1.368559E-4   1.489835E+0   9.148983E+1   
2.168546E+3   1.199599E+2   1.199599E+2   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   9.796200E-2   -1.161195E-1   1.361921E-4   3.459940E-6   -3.459940E-6   1.361921E-4   1.362361E-4   1.455278E+0   9.145528E+1   
2.190874E+3   1.199889E+2   1.199889E+2   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   9.765828E-2   -1.165681E-1   1.362965E-4   3.977831E-6   -3.977831E-6   1.362965E-4   1.363545E-4   1.671710E+0   9.167171E+1   
2.213105E+3   1.200383E+2   1.200383E+2   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   9.695998E-2   -1.166666E-1   1.359289E-4   4.558686E-6   -4.558686E-6   1.359289E-4   1.360053E-4   1.920825E+0   9.192083E+1   
2.235339E+3   1.200711E+2   1.200711E+2   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.400000E+1   -3.400000E+1   9.804207E-2   -1.170706E-1   1.368610E-4   4.022493E-6   -4.022493E-6   1.368610E-4   1.369201E-4   1.683500E+0   9.168350E+1   
2.257621E+3   1.200724E+2   1.200724E+2   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   9.782180E-2   -1.172446E-1   1.368382E-4   4.299145E-6   -4.299145E-6   1.368382E-4   1.369057E-4   1.799512E+0   9.179951E+1   
2.279838E+3   1.201002E+2   1.201002E+2   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   9.860444E-2   -1.160278E-1   1.365296E-4   2.924810E-6   -2.924810E-6   1.365296E-4   1.365609E-4   1.227233E+0   9.122723E+1   
2.302090E+3   1.200206E+2   1.200206E+2   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   9.932540E-2   -1.164527E-1   1.372520E-4   2.669365E-6   -2.669365E-6   1.372520E-4   1.372780E-4   1.114184E+0   9.111418E+1   
2.324328E+3   1.200413E+2   1.200413E+2   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   9.842714E-2   -1.172811E-1   1.372362E-4   3.875283E-6   -3.875283E-6   1.372362E-4   1.372909E-4   1.617492E+0   9.161749E+1   
2.346592E+3   1.200419E+2   1.200419E+2   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   9.815282E-2   -1.167724E-1   1.367353E-4   3.745629E-6   -3.745629E-6   1.367353E-4   1.367866E-4   1.569127E+0   9.156913E+1   
2.368831E+3   1.200326E+2   1.200326E+2   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   9.805311E-2   -1.167114E-1   1.366339E-4   3.779465E-6   -3.779465E-6   1.366339E-4   1.366861E-4   1.584469E+0   9.158447E+1   
2.391022E+3   1.200901E+2   1.200901E+2   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   9.800465E-2   -1.165150E-1   1.364761E-4   3.686936E-6   -3.686936E-6   1.364761E-4   1.365258E-4   1.547484E+0   9.154748E+1   
2.424387E+3   1.200059E+2   1.200059E+2   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   9.989943E-2   -1.184742E-1   1.389235E-4   3.566355E-6   -3.566355E-6   1.389235E-4   1.389692E-4   1.470538E+0   9.147054E+1   
2.446046E+3   1.200680E+2   1.200680E+2   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   1.015564E-1   -1.197284E-1   1.407647E-4   3.160742E-6   -3.160742E-6   1.407647E-4   1.408002E-4   1.286307E+0   9.128631E+1   
2.467765E+3   1.200600E+2   1.200600E+2   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   1.020494E-1   -1.218241E-1   1.424344E-4   4.166205E-6   -4.166205E-6   1.424344E-4   1.424954E-4   1.675423E+0   9.167542E+1   
2.489496E+3   1.200919E+2   1.200919E+2   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   1.035450E-1   -1.230169E-1   1.441360E-4   3.839824E-6   -3.839824E-6   1.441360E-4   1.441871E-4   1.526015E+0   9.152602E+1   
2.511232E+3   1.200094E+2   1.200094E+2   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   1.042341E-1   -1.250491E-1   1.458855E-4   4.658760E-6   -4.658760E-6   1.458855E-4   1.459599E-4   1.829082E+0   9.182908E+1   
2.532958E+3   1.199976E+2   1.199976E+2   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   1.069348E-1   -1.270457E-1   1.488556E-4   3.966569E-6   -3.966569E-6   1.488556E-4   1.489084E-4   1.526405E+0   9.152640E+1   
2.554722E+3   1.201141E+2   1.201141E+2   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   1.063795E-1   -1.281406E-1   1.492254E-4   5.093120E-6   -5.093120E-6   1.492254E-4   1.493123E-4   1.954768E+0   9.195477E+1   
2.576433E+3   1.201013E+2   1.201013E+2   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   1.079015E-1   -1.291607E-1   1.508307E-4   4.634309E-6   -4.634309E-6   1.508307E-4   1.509019E-4   1.759873E+0   9.175987E+1   
2.598170E+3   1.199769E+2   1.199769E+2   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   1.091977E-1   -1.316003E-1   1.532210E-4   5.270550E-6   -5.270550E-6   1.532210E-4   1.533116E-4   1.970104E+0   9.197010E+1   
2.619902E+3   1.200671E+2   1.200671E+2   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   1.099947E-1   -1.340853E-1   1.553322E-4   6.305668E-6   -6.305668E-6   1.553322E-4   1.554602E-4   2.324629E+0   9.232463E+1   
2.641629E+3   1.200243E+2   1.200243E+2   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   1.111234E-1   -1.345127E-1   1.563084E-4   5.750247E-6   -5.750247E-6   1.563084E-4   1.564141E-4   2.106838E+0   9.210684E+1   
2.663353E+3   1.200258E+2   1.200258E+2   -6.510000E+2   -6.510000E+2   9.000000E+1   -6.500000E+2   -6.500000E+2   1.125552E-1   -1.370812E-1   1.588664E-4   6.370441E-6   -6.370441E-6   1.588664E-4   1.589941E-4   2.296293E+0   9.229629E+1   
2.684981E+3   1.199829E+2   1.199829E+2   -7.010000E+2   -7.010000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   1.134793E-1   -1.388529E-1   1.605916E-4   6.845271E-6   -6.845271E-6   1.605916E-4   1.607374E-4   2.440774E+0   9.244077E+1   
2.706662E+3   1.200478E+2   1.200478E+2   -7.510000E+2   -7.510000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   1.135885E-1   -1.413526E-1   1.622872E-4   8.398755E-6   -8.398755E-6   1.622872E-4   1.625044E-4   2.962552E+0   9.296255E+1   
2.728454E+3   1.200107E+2   1.200107E+2   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   1.148952E-1   -1.421104E-1   1.635886E-4   7.927743E-6   -7.927743E-6   1.635886E-4   1.637805E-4   2.774467E+0   9.277447E+1   
2.750129E+3   1.200185E+2   1.200185E+2   -8.510000E+2   -8.510000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   1.165659E-1   -1.446101E-1   1.662496E-4   8.326248E-6   -8.326248E-6   1.662496E-4   1.664579E-4   2.867139E+0   9.286714E+1   
2.771855E+3   1.200188E+2   1.200188E+2   -9.000000E+2   -9.000000E+2   9.000000E+1   -9.000000E+2   -9.000000E+2   1.196170E-1   -1.449074E-1   1.683295E-4   6.263929E-6   -6.263929E-6   1.683295E-4   1.684460E-4   2.131125E+0   9.213113E+1   
2.793487E+3   1.200491E+2   1.200491E+2   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.490000E+2   -9.490000E+2   1.221449E-1   -1.470749E-1   1.713041E-4   5.811235E-6   -5.811235E-6   1.713041E-4   1.714026E-4   1.942929E+0   9.194293E+1   
2.815189E+3   1.201014E+2   1.201014E+2   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   1.208657E-1   -1.490378E-1   1.717915E-4   8.040691E-6   -8.040691E-6   1.717915E-4   1.719796E-4   2.679770E+0   9.267977E+1   
2.836957E+3   1.200124E+2   1.200124E+2   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   1.217016E-1   -1.506113E-1   1.733332E-4   8.451111E-6   -8.451111E-6   1.733332E-4   1.735391E-4   2.791328E+0   9.279133E+1   
2.858826E+3   1.200640E+2   1.200640E+2   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   1.227702E-1   -1.523600E-1   1.751328E-4   8.804035E-6   -8.804035E-6   1.751328E-4   1.753539E-4   2.877873E+0   9.287787E+1   
2.880636E+3   1.200301E+2   1.200301E+2   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   1.235320E-1   -1.551801E-1   1.774404E-4   1.008426E-5   -1.008426E-5   1.774404E-4   1.777267E-4   3.252726E+0   9.325273E+1   
2.903020E+3   1.200247E+2   1.200247E+2   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   1.264769E-1   -1.559526E-1   1.797642E-4   8.411175E-6   -8.411175E-6   1.797642E-4   1.799609E-4   2.678918E+0   9.267892E+1   
2.924893E+3   1.200224E+2   1.200224E+2   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   1.270561E-1   -1.578418E-1   1.813527E-4   9.217893E-6   -9.217893E-6   1.813527E-4   1.815868E-4   2.909757E+0   9.290976E+1   
2.946768E+3   1.200755E+2   1.200755E+2   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   1.288306E-1   -1.599470E-1   1.838209E-4   9.281726E-6   -9.281726E-6   1.838209E-4   1.840551E-4   2.890599E+0   9.289060E+1   
2.969382E+3   1.200945E+2   1.200945E+2   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   1.292337E-1   -1.614727E-1   1.850638E-4   9.981021E-6   -9.981021E-6   1.850638E-4   1.853327E-4   3.087135E+0   9.308713E+1   
2.991305E+3   1.200026E+2   1.200026E+2   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   1.305238E-1   -1.626039E-1   1.865981E-4   9.766377E-6   -9.766377E-6   1.865981E-4   1.868535E-4   2.996077E+0   9.299608E+1   
3.013113E+3   1.200005E+2   1.200005E+2   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   1.323661E-1   -1.654635E-1   1.895995E-4   1.027328E-5   -1.027328E-5   1.895995E-4   1.898776E-4   3.101487E+0   9.310149E+1   
3.035947E+3   1.200866E+2   1.200866E+2   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   1.326330E-1   -1.669459E-1   1.907300E-4   1.104502E-5   -1.104502E-5   1.907300E-4   1.910495E-4   3.314250E+0   9.331425E+1   
3.058031E+3   1.200377E+2   1.200377E+2   -1.550000E+3   -1.550000E+3   9.000000E+1   -1.548000E+3   -1.548000E+3   1.347578E-1   -1.692668E-1   1.935552E-4   1.099077E-5   -1.099077E-5   1.935552E-4   1.938670E-4   3.249972E+0   9.324997E+1   
3.080163E+3   1.200084E+2   1.200084E+2   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   1.362718E-1   -1.712931E-1   1.958110E-4   1.119573E-5   -1.119573E-5   1.958110E-4   1.961308E-4   3.272392E+0   9.327239E+1   
3.102582E+3   1.199658E+2   1.199658E+2   -1.650000E+3   -1.650000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   1.345016E-1   -1.724752E-1   1.954865E-4   1.327783E-5   -1.327783E-5   1.954865E-4   1.959369E-4   3.885674E+0   9.388567E+1   
3.124711E+3   1.200270E+2   1.200270E+2   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   1.387372E-1   -1.737582E-1   1.989407E-4   1.098386E-5   -1.098386E-5   1.989407E-4   1.992437E-4   3.160189E+0   9.316019E+1   
3.146847E+3   1.199950E+2   1.199950E+2   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   1.382457E-1   -1.744970E-1   1.991180E-4   1.183034E-5   -1.183034E-5   1.991180E-4   1.994691E-4   3.400158E+0   9.340016E+1   
3.170005E+3   1.199862E+2   1.199862E+2   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.799000E+3   -1.799000E+3   1.394956E-1   -1.757702E-1   2.007200E-4   1.173828E-5   -1.173828E-5   2.007200E-4   2.010629E-4   3.346895E+0   9.334689E+1   
3.192147E+3   1.200213E+2   1.200213E+2   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.848000E+3   -1.848000E+3   1.403540E-1   -1.771286E-1   2.021354E-4   1.199151E-5   -1.199151E-5   2.021354E-4   2.024908E-4   3.395043E+0   9.339504E+1   
3.214279E+3   1.200391E+2   1.200391E+2   -1.900000E+3   -1.900000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   1.414296E-1   -1.789948E-1   2.040159E-4   1.241603E-5   -1.241603E-5   2.040159E-4   2.043933E-4   3.482620E+0   9.348262E+1   
3.237463E+3   1.200560E+2   1.200560E+2   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   1.421481E-1   -1.807773E-1   2.056210E-4   1.304992E-5   -1.304992E-5   2.056210E-4   2.060347E-4   3.631458E+0   9.363146E+1   
3.259830E+3   1.200186E+2   1.200186E+2   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   1.431814E-1   -1.818738E-1   2.069740E-4   1.300253E-5   -1.300253E-5   2.069740E-4   2.073820E-4   3.594716E+0   9.359472E+1   
3.296870E+3   1.199926E+2   1.199926E+2   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.544441E-1   -1.994795E-1   2.254034E-4   1.618242E-5   -1.618242E-5   2.254034E-4   2.259836E-4   4.106399E+0   9.410640E+1   
3.322966E+3   1.200675E+2   1.200675E+2   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.641933E-1   -2.162788E-1   2.423721E-4   1.995452E-5   -1.995452E-5   2.423721E-4   2.431922E-4   4.706551E+0   9.470655E+1   
3.348139E+3   1.200733E+2   1.200733E+2   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.760174E-1   -2.352316E-1   2.620260E-4   2.359981E-5   -2.359981E-5   2.620260E-4   2.630867E-4   5.146553E+0   9.514655E+1   
3.373738E+3   1.200128E+2   1.200128E+2   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   1.883232E-1   -2.509515E-1   2.798723E-4   2.477526E-5   -2.477526E-5   2.798723E-4   2.809667E-4   5.058834E+0   9.505883E+1   
3.399400E+3   1.200463E+2   1.200463E+2   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   1.911754E-1   -2.599336E-1   2.874855E-4   2.853802E-5   -2.853802E-5   2.874855E-4   2.888985E-4   5.669046E+0   9.566905E+1   
3.424131E+3   1.200524E+2   1.200524E+2   -5.000000E+3   -5.000000E+3   9.000000E+1   -5.000000E+3   -5.000000E+3   1.851931E-1   -2.568243E-1   2.817620E-4   3.092989E-5   -3.092989E-5   2.817620E-4   2.834546E-4   6.264454E+0   9.626445E+1   
3.449276E+3   1.200733E+2   1.200733E+2   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   1.763006E-1   -2.440819E-1   2.679652E-4   2.917648E-5   -2.917648E-5   2.679652E-4   2.695489E-4   6.213976E+0   9.621398E+1   
3.475457E+3   1.200440E+2   1.200440E+2   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   1.589533E-1   -2.243082E-1   2.443619E-4   2.907956E-5   -2.907956E-5   2.443619E-4   2.460861E-4   6.786398E+0   9.678640E+1   
3.500153E+3   1.200639E+2   1.200639E+2   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.474624E-1   -2.128170E-1   2.297736E-4   3.006595E-5   -3.006595E-5   2.297736E-4   2.317323E-4   7.454816E+0   9.745482E+1   
3.524886E+3   1.201004E+2   1.201004E+2   -7.001000E+3   -7.001000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.428562E-1   -2.079862E-1   2.237796E-4   3.031463E-5   -3.031463E-5   2.237796E-4   2.258236E-4   7.714694E+0   9.771469E+1   
3.549661E+3   1.200380E+2   1.200380E+2   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.458837E-1   -2.157601E-1   2.307143E-4   3.315775E-5   -3.315775E-5   2.307143E-4   2.330848E-4   8.178421E+0   9.817842E+1   
3.574892E+3   1.200107E+2   1.200107E+2   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.490396E-1   -2.230359E-1   2.374042E-4   3.558026E-5   -3.558026E-5   2.374042E-4   2.400557E-4   8.523597E+0   9.852360E+1   
3.600151E+3   1.200412E+2   1.200412E+2   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.610904E-1   -2.387830E-1   2.551105E-4   3.696209E-5   -3.696209E-5   2.551105E-4   2.577742E-4   8.244024E+0   9.824402E+1   
3.625801E+3   1.200654E+2   1.200654E+2   -9.000000E+3   -9.000000E+3   9.000000E+1   -9.000000E+3   -9.000000E+3   1.749498E-1   -2.546445E-1   2.740094E-4   3.708108E-5   -3.708108E-5   2.740094E-4   2.765071E-4   7.706890E+0   9.770689E+1   
3.650969E+3   1.200194E+2   1.200194E+2   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.847348E-1   -2.718399E-1   2.912581E-4   4.108565E-5   -4.108565E-5   2.912581E-4   2.941417E-4   8.029319E+0   9.802932E+1   
3.676145E+3   1.200307E+2   1.200307E+2   -1.000000E+4   -1.000000E+4   9.000000E+1   -9.999000E+3   -9.999000E+3   2.040120E-1   -2.944443E-1   3.178983E-4   4.160575E-5   -4.160575E-5   3.178983E-4   3.206093E-4   7.456351E+0   9.745635E+1   
3.712643E+3   1.200266E+2   1.200266E+2   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.832165E-1   -2.670037E-1   2.871697E-4   3.904687E-5   -3.904687E-5   2.871697E-4   2.898121E-4   7.743104E+0   9.774310E+1   
3.737274E+3   1.200378E+2   1.200378E+2   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.775459E-1   -2.552859E-1   2.760322E-4   3.558028E-5   -3.558028E-5   2.760322E-4   2.783158E-4   7.344872E+0   9.734487E+1   
3.761518E+3   1.199737E+2   1.199737E+2   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.560661E-1   -2.307610E-1   2.467796E-4   3.543369E-5   -3.543369E-5   2.467796E-4   2.493104E-4   8.170933E+0   9.817093E+1   
3.786174E+3   1.200079E+2   1.200079E+2   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.471163E-1   -2.149461E-1   2.309463E-4   3.171389E-5   -3.171389E-5   2.309463E-4   2.331137E-4   7.819036E+0   9.781904E+1   
3.810966E+3   1.200391E+2   1.200391E+2   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.345851E-1   -1.966693E-1   2.112954E-4   2.903350E-5   -2.903350E-5   2.112954E-4   2.132808E-4   7.823854E+0   9.782385E+1   
3.836107E+3   1.200174E+2   1.200174E+2   -7.000000E+3   -7.000000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.148807E-1   -1.746939E-1   1.848009E-4   2.924061E-5   -2.924061E-5   1.848009E-4   1.871000E-4   8.991233E+0   9.899123E+1   
3.860819E+3   1.201209E+2   1.201209E+2   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.013245E-1   -1.559480E-1   1.642108E-4   2.701168E-5   -2.701168E-5   1.642108E-4   1.664176E-4   9.341155E+0   9.934116E+1   
3.885006E+3   1.199757E+2   1.199757E+2   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   8.762249E-2   -1.365200E-1   1.430864E-4   2.444463E-5   -2.444463E-5   1.430864E-4   1.451594E-4   9.694719E+0   9.969472E+1   
3.909657E+3   1.200908E+2   1.200908E+2   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   6.951248E-2   -1.146700E-1   1.176592E-4   2.355438E-5   -2.355438E-5   1.176592E-4   1.199937E-4   1.132049E+1   1.013205E+2   
3.934812E+3   1.200641E+2   1.200641E+2   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   5.916315E-2   -9.630893E-2   9.930241E-5   1.920516E-5   -1.920516E-5   9.930241E-5   1.011425E-4   1.094591E+1   1.009459E+2   
3.959549E+3   1.200152E+2   1.200152E+2   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   4.485946E-2   -7.718509E-2   7.800404E-5   1.728199E-5   -1.728199E-5   7.800404E-5   7.989554E-5   1.249223E+1   1.024922E+2   
3.984180E+3   1.200859E+2   1.200859E+2   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   3.463399E-2   -5.951903E-2   6.017647E-5   1.329549E-5   -1.329549E-5   6.017647E-5   6.162773E-5   1.245887E+1   1.024589E+2   
4.008881E+3   1.200535E+2   1.200535E+2   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   2.085894E-2   -4.075389E-2   3.943855E-5   1.121583E-5   -1.121583E-5   3.943855E-5   4.100237E-5   1.587509E+1   1.058751E+2   
4.033046E+3   1.199994E+2   1.199994E+2   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   8.179441E-3   -2.260490E-2   1.977925E-5   8.728679E-6   -8.728679E-6   1.977925E-5   2.161963E-5   2.381210E+1   1.138121E+2   
4.058196E+3   1.200696E+2   1.200696E+2   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   -3.803943E-3   -3.951511E-3   2.218016E-7   5.396901E-6   -5.396901E-6   2.218016E-7   5.401457E-6   8.764658E+1   1.776466E+2   
4.082868E+3   1.199873E+2   1.199873E+2   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   -1.696327E-2   1.459390E-2   -1.999234E-5   3.005479E-6   -3.005479E-6   -1.999234E-5   2.021698E-5   1.714507E+2   2.614507E+2   
4.116553E+3   1.199901E+2   1.199901E+2   -1.950000E+3   -1.950000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   -1.594348E-2   1.648375E-2   -2.059270E-5   1.015688E-6   -1.015688E-6   -2.059270E-5   2.061773E-5   1.771763E+2   2.671763E+2   
4.138561E+3   1.200453E+2   1.200453E+2   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.899000E+3   -1.899000E+3   -1.683748E-2   1.811374E-2   -2.220701E-5   6.112727E-7   -6.112727E-7   -2.220701E-5   2.221542E-5   1.784233E+2   2.684233E+2   
4.160589E+3   1.200756E+2   1.200756E+2   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.849000E+3   -1.849000E+3   -1.929121E-2   1.865155E-2   -2.407428E-5   2.074520E-6   -2.074520E-6   -2.407428E-5   2.416350E-5   1.750749E+2   2.650749E+2   
4.182475E+3   1.200642E+2   1.200642E+2   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.799000E+3   -1.799000E+3   -1.794439E-2   2.033492E-2   -2.433798E-5   -2.217074E-8   2.217074E-8   -2.433798E-5   2.433799E-5   -1.799478E+2   -8.994781E+1   
4.204504E+3   1.199921E+2   1.199921E+2   -1.750000E+3   -1.750000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   -2.080708E-2   2.271535E-2   -2.765818E-5   5.389071E-7   -5.389071E-7   -2.765818E-5   2.766343E-5   1.788838E+2   2.688838E+2   
4.226590E+3   1.200384E+2   1.200384E+2   -1.700000E+3   -1.700000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   -2.036714E-2   2.594347E-2   -2.948862E-5   -1.896935E-6   1.896935E-6   -2.948862E-5   2.954957E-5   -1.763194E+2   -8.631937E+1   
4.248427E+3   1.201043E+2   1.201043E+2   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   -2.157745E-2   2.633095E-2   -3.048925E-5   -1.255081E-6   1.255081E-6   -3.048925E-5   3.051507E-5   -1.776428E+2   -8.764277E+1   
4.270247E+3   1.200275E+2   1.200275E+2   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.599000E+3   -1.599000E+3   -2.279634E-2   2.743939E-2   -3.196475E-5   -1.078217E-6   1.078217E-6   -3.196475E-5   3.198293E-5   -1.780681E+2   -8.806806E+1   
4.292361E+3   1.200388E+2   1.200388E+2   -1.550000E+3   -1.550000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   -2.415177E-2   3.021494E-2   -3.461043E-5   -1.890274E-6   1.890274E-6   -3.461043E-5   3.466201E-5   -1.768739E+2   -8.687386E+1   
4.314168E+3   1.200315E+2   1.200315E+2   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   -2.572225E-2   3.045548E-2   -3.573803E-5   -8.859559E-7   8.859559E-7   -3.573803E-5   3.574901E-5   -1.785799E+2   -8.857991E+1   
4.336291E+3   1.200124E+2   1.200124E+2   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   -2.581492E-2   3.326049E-2   -3.762220E-5   -2.651247E-6   2.651247E-6   -3.762220E-5   3.771550E-5   -1.759690E+2   -8.596901E+1   
4.358323E+3   1.200435E+2   1.200435E+2   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   -2.663344E-2   3.465179E-2   -3.903438E-5   -2.955439E-6   2.955439E-6   -3.903438E-5   3.914611E-5   -1.756702E+2   -8.567018E+1   
4.380440E+3   1.200589E+2   1.200589E+2   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   -2.869541E-2   3.737119E-2   -4.208031E-5   -3.208210E-6   3.208210E-6   -4.208031E-5   4.220243E-5   -1.756402E+2   -8.564019E+1   
4.402432E+3   1.199711E+2   1.199711E+2   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.300000E+3   -1.300000E+3   -3.026037E-2   3.782370E-2   -4.334255E-5   -2.346560E-6   2.346560E-6   -4.334255E-5   4.340602E-5   -1.769010E+2   -8.690104E+1   
4.424552E+3   1.200586E+2   1.200586E+2   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   -3.047358E-2   3.828238E-2   -4.377310E-5   -2.488732E-6   2.488732E-6   -4.377310E-5   4.384379E-5   -1.767459E+2   -8.674593E+1   
4.446638E+3   1.200055E+2   1.200055E+2   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   -3.226431E-2   4.227252E-2   -4.747895E-5   -3.772888E-6   3.772888E-6   -4.747895E-5   4.762862E-5   -1.754566E+2   -8.545657E+1   
4.468642E+3   1.200574E+2   1.200574E+2   -1.151000E+3   -1.151000E+3   9.000000E+1   -1.150000E+3   -1.150000E+3   -3.422933E-2   4.392429E-2   -4.976960E-5   -3.399384E-6   3.399384E-6   -4.976960E-5   4.988556E-5   -1.760926E+2   -8.609263E+1   
4.490717E+3   1.200215E+2   1.200215E+2   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.100000E+3   -1.100000E+3   -3.571207E-2   4.425106E-2   -5.089912E-5   -2.516339E-6   2.516339E-6   -5.089912E-5   5.096128E-5   -1.771697E+2   -8.716973E+1   
4.512770E+3   1.200479E+2   1.200479E+2   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.050000E+3   -1.050000E+3   -3.689506E-2   4.626182E-2   -5.294009E-5   -2.955941E-6   2.955941E-6   -5.294009E-5   5.302255E-5   -1.768042E+2   -8.680418E+1   
4.534848E+3   1.200164E+2   1.200164E+2   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   -3.736567E-2   4.903804E-2   -5.503916E-5   -4.422876E-6   4.422876E-6   -5.503916E-5   5.521658E-5   -1.754057E+2   -8.540566E+1   
4.556817E+3   1.200219E+2   1.200219E+2   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   -4.020382E-2   4.991947E-2   -5.736790E-5   -2.899944E-6   2.899944E-6   -5.736790E-5   5.744115E-5   -1.771062E+2   -8.710617E+1   
4.578412E+3   1.200457E+2   1.200457E+2   -9.000000E+2   -9.000000E+2   9.000000E+1   -9.000000E+2   -9.000000E+2   -4.060388E-2   5.190506E-2   -5.890843E-5   -3.902173E-6   3.902173E-6   -5.890843E-5   5.903753E-5   -1.762102E+2   -8.621019E+1   
4.600292E+3   1.200037E+2   1.200037E+2   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   -3.996880E-2   5.342981E-2   -5.950885E-5   -5.368733E-6   5.368733E-6   -5.950885E-5   5.975054E-5   -1.748449E+2   -8.484488E+1   
4.621918E+3   1.200124E+2   1.200124E+2   -8.000000E+2   -8.000000E+2   9.000000E+1   -8.000000E+2   -8.000000E+2   -4.222344E-2   5.526750E-2   -6.209964E-5   -4.902567E-6   4.902567E-6   -6.209964E-5   6.229286E-5   -1.754860E+2   -8.548604E+1   
4.643642E+3   1.200040E+2   1.200040E+2   -7.500000E+2   -7.500000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   -4.470572E-2   5.708617E-2   -6.481879E-5   -4.255583E-6   4.255583E-6   -6.481879E-5   6.495833E-5   -1.762437E+2   -8.624372E+1   
4.665576E+3   1.200593E+2   1.200593E+2   -7.010000E+2   -7.010000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   -4.365218E-2   5.823911E-2   -6.491833E-5   -5.788574E-6   5.788574E-6   -6.491833E-5   6.517590E-5   -1.749046E+2   -8.490458E+1   
4.687556E+3   1.200744E+2   1.200744E+2   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.500000E+2   -6.500000E+2   -4.487567E-2   6.074158E-2   -6.730459E-5   -6.519690E-6   6.519690E-6   -6.730459E-5   6.761963E-5   -1.744671E+2   -8.446711E+1   
4.709178E+3   1.200330E+2   1.200330E+2   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   -4.754147E-2   6.264003E-2   -7.018915E-5   -5.789136E-6   5.789136E-6   -7.018915E-5   7.042748E-5   -1.752850E+2   -8.528497E+1   
4.730817E+3   1.200572E+2   1.200572E+2   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   -4.875700E-2   6.392856E-2   -7.177985E-5   -5.732495E-6   5.732495E-6   -7.177985E-5   7.200839E-5   -1.754339E+2   -8.543393E+1   
4.752511E+3   1.200162E+2   1.200162E+2   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   -4.785226E-2   6.457834E-2   -7.164369E-5   -6.826475E-6   6.826475E-6   -7.164369E-5   7.196818E-5   -1.745571E+2   -8.455708E+1   
4.774181E+3   1.200652E+2   1.200652E+2   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   -5.139732E-2   6.670964E-2   -7.522351E-5   -5.597824E-6   5.597824E-6   -7.522351E-5   7.543150E-5   -1.757441E+2   -8.574413E+1   
4.795813E+3   1.200693E+2   1.200693E+2   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   -5.167466E-2   6.759045E-2   -7.596863E-5   -5.968544E-6   5.968544E-6   -7.596863E-5   7.620273E-5   -1.755077E+2   -8.550773E+1   
4.817518E+3   1.199870E+2   1.199870E+2   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   -5.136755E-2   7.086483E-2   -7.791133E-5   -8.336391E-6   8.336391E-6   -7.791133E-5   7.835605E-5   -1.738927E+2   -8.389268E+1   
4.839230E+3   1.200308E+2   1.200308E+2   -3.000000E+2   -3.000000E+2   9.000000E+1   -3.000000E+2   -3.000000E+2   -5.294723E-2   7.099216E-2   -7.897090E-5   -7.251253E-6   7.251253E-6   -7.897090E-5   7.930311E-5   -1.747537E+2   -8.475371E+1   
4.860873E+3   1.199889E+2   1.199889E+2   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   -5.248735E-2   7.284610E-2   -7.989403E-5   -8.803445E-6   8.803445E-6   -7.989403E-5   8.037759E-5   -1.737120E+2   -8.371200E+1   
4.882595E+3   1.199922E+2   1.199922E+2   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   -5.656708E-2   7.387600E-2   -8.308707E-5   -6.459270E-6   6.459270E-6   -8.308707E-5   8.333777E-5   -1.755547E+2   -8.555471E+1   
4.904276E+3   1.199716E+2   1.199716E+2   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   -5.683245E-2   7.603214E-2   -8.465541E-5   -7.672621E-6   7.672621E-6   -8.465541E-5   8.500240E-5   -1.748212E+2   -8.482123E+1   
4.925956E+3   1.200776E+2   1.200776E+2   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   -5.705182E-2   7.779191E-2   -8.593715E-5   -8.660853E-6   8.660853E-6   -8.593715E-5   8.637248E-5   -1.742451E+2   -8.424509E+1   
4.947474E+3   1.199950E+2   1.199950E+2   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   -5.887323E-2   7.830793E-2   -8.739931E-5   -7.651041E-6   7.651041E-6   -8.739931E-5   8.773356E-5   -1.749970E+2   -8.499701E+1   
4.980509E+3   1.200342E+2   1.200342E+2   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   -5.925183E-2   7.937802E-2   -8.833031E-5   -8.070614E-6   8.070614E-6   -8.833031E-5   8.869824E-5   -1.747795E+2   -8.477946E+1   
5.002779E+3   1.200264E+2   1.200264E+2   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   -5.861186E-2   8.030883E-2   -8.854088E-5   -9.152491E-6   9.152491E-6   -8.854088E-5   8.901268E-5   -1.740983E+2   -8.409828E+1   
5.024974E+3   1.200372E+2   1.200372E+2   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   -5.788291E-2   7.927248E-2   -8.741525E-5   -9.014108E-6   9.014108E-6   -8.741525E-5   8.787878E-5   -1.741126E+2   -8.411257E+1   
5.047255E+3   1.200120E+2   1.200120E+2   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   -5.922422E-2   7.844261E-2   -8.770402E-5   -7.479488E-6   7.479488E-6   -8.770402E-5   8.802237E-5   -1.751256E+2   -8.512555E+1   
5.069487E+3   1.200460E+2   1.200460E+2   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   -5.811116E-2   7.897366E-2   -8.736175E-5   -8.649930E-6   8.649930E-6   -8.736175E-5   8.778893E-5   -1.743454E+2   -8.434542E+1   
5.091741E+3   1.199817E+2   1.199817E+2   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   -5.755680E-2   7.920498E-2   -8.716967E-5   -9.211181E-6   9.211181E-6   -8.716967E-5   8.765499E-5   -1.739680E+2   -8.396796E+1   
5.114016E+3   1.199349E+2   1.199349E+2   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   -5.857901E-2   7.908626E-2   -8.772433E-5   -8.377507E-6   8.377507E-6   -8.772433E-5   8.812344E-5   -1.745449E+2   -8.454490E+1   
5.136269E+3   1.200349E+2   1.200349E+2   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   -5.934938E-2   7.954462E-2   -8.849913E-5   -8.107383E-6   8.107383E-6   -8.849913E-5   8.886971E-5   -1.747658E+2   -8.476576E+1   
5.158523E+3   1.200370E+2   1.200370E+2   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   -5.844188E-2   7.991430E-2   -8.817884E-5   -9.020279E-6   9.020279E-6   -8.817884E-5   8.863901E-5   -1.741592E+2   -8.415923E+1   
5.180762E+3   1.200699E+2   1.200699E+2   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   -5.781696E-2   7.978790E-2   -8.771016E-5   -9.399861E-6   9.399861E-6   -8.771016E-5   8.821241E-5   -1.738830E+2   -8.388298E+1   
5.202994E+3   1.200644E+2   1.200644E+2   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   -5.925184E-2   7.973207E-2   -8.856091E-5   -8.302077E-6   8.302077E-6   -8.856091E-5   8.894919E-5   -1.746445E+2   -8.464450E+1   
5.225279E+3   1.199790E+2   1.199790E+2   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   -5.864344E-2   8.031865E-2   -8.856680E-5   -9.135551E-6   9.135551E-6   -8.856680E-5   8.903672E-5   -1.741108E+2   -8.411084E+1   
5.247587E+3   1.200568E+2   1.200568E+2   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   -5.858333E-2   7.982287E-2   -8.820675E-5   -8.855885E-6   8.855885E-6   -8.820675E-5   8.865020E-5   -1.742668E+2   -8.426676E+1   
5.269776E+3   1.199774E+2   1.199774E+2   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   -5.834310E-2   8.041744E-2   -8.844546E-5   -9.422280E-6   9.422280E-6   -8.844546E-5   8.894594E-5   -1.739191E+2   -8.391910E+1   
5.292071E+3   1.199983E+2   1.199983E+2   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   -5.846797E-2   7.953295E-2   -8.794660E-5   -8.751670E-6   8.751670E-6   -8.794660E-5   8.838097E-5   -1.743171E+2   -8.431714E+1   
5.314313E+3   1.200975E+2   1.200975E+2   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   -5.799612E-2   7.988854E-2   -8.788647E-5   -9.333133E-6   9.333133E-6   -8.788647E-5   8.838065E-5   -1.739382E+2   -8.393818E+1   
5.336588E+3   1.200388E+2   1.200388E+2   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   -5.870634E-2   7.863436E-2   -8.750873E-5   -7.987889E-6   7.987889E-6   -8.750873E-5   8.787255E-5   -1.747844E+2   -8.478443E+1   
5.358793E+3   1.200319E+2   1.200319E+2   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   -5.874744E-2   8.039105E-2   -8.867825E-5   -9.105961E-6   9.105961E-6   -8.867825E-5   8.914455E-5   -1.741371E+2   -8.413711E+1   
5.381037E+3   1.200358E+2   1.200358E+2   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   -5.805319E-2   8.062145E-2   -8.839909E-5   -9.770085E-6   9.770085E-6   -8.839909E-5   8.893736E-5   -1.736931E+2   -8.369313E+1   
5.403182E+3   1.199969E+2   1.199969E+2   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   -5.735278E-2   8.088468E-2   -8.813750E-5   -1.046022E-5   1.046022E-5   -8.813750E-5   8.875605E-5   -1.732318E+2   -8.323175E+1   
5.425264E+3   1.200378E+2   1.200378E+2   -8.000000E+0   -8.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   -5.868304E-2   7.992963E-2   -8.833792E-5   -8.851931E-6   8.851931E-6   -8.833792E-5   8.878032E-5   -1.742778E+2   -8.427776E+1   
5.447286E+3   1.200381E+2   1.200381E+2   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   -5.922911E-2   7.983944E-2   -8.861679E-5   -8.389079E-6   8.389079E-6   -8.861679E-5   8.901299E-5   -1.745921E+2   -8.459210E+1   
5.469378E+3   1.200566E+2   1.200566E+2   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   -5.812497E-2   8.054504E-2   -8.839371E-5   -9.667045E-6   9.667045E-6   -8.839371E-5   8.892075E-5   -1.737587E+2   -8.375874E+1   
5.491475E+3   1.199611E+2   1.199611E+2   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   -5.892571E-2   8.086627E-2   -8.909797E-5   -9.284801E-6   9.284801E-6   -8.909797E-5   8.958045E-5   -1.740507E+2   -8.405074E+1   
5.513518E+3   1.199908E+2   1.199908E+2   0.000000E+0   0.000000E+0   9.000000E+1   0.000000E+0   0.000000E+0   -5.968593E-2   7.953570E-2   -8.870139E-5   -7.852627E-6   7.852627E-6   -8.870139E-5   8.904831E-5   -1.749409E+2   -8.494086E+1   
5.535509E+3   1.199537E+2   1.199537E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   -5.815012E-2   8.017076E-2   -8.816549E-5   -9.403738E-6   9.403738E-6   -8.816549E-5   8.866557E-5   -1.739118E+2   -8.391184E+1   
5.557052E+3   1.200224E+2   1.200224E+2   3.000000E+0   3.000000E+0   9.000000E+1   3.000000E+0   3.000000E+0   -6.021883E-2   8.066317E-2   -8.976517E-5   -8.195583E-6   8.195583E-6   -8.976517E-5   9.013852E-5   -1.747833E+2   -8.478334E+1   
5.578730E+3   1.199667E+2   1.199667E+2   5.000000E+0   5.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   -5.881250E-2   8.035302E-2   -8.869370E-5   -9.032983E-6   9.032983E-6   -8.869370E-5   8.915250E-5   -1.741848E+2   -8.418478E+1   
5.600453E+3   1.199839E+2   1.199839E+2   7.000000E+0   7.000000E+0   9.000000E+1   8.000000E+0   8.000000E+0   -5.868888E-2   7.999192E-2   -8.838210E-5   -8.888337E-6   8.888337E-6   -8.838210E-5   8.882791E-5   -1.742572E+2   -8.425723E+1   
5.622133E+3   1.199493E+2   1.199493E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   -5.786913E-2   8.142309E-2   -8.880740E-5   -1.043031E-5   1.043031E-5   -8.880740E-5   8.941781E-5   -1.733014E+2   -8.330137E+1   
5.643966E+3   1.200121E+2   1.200121E+2   1.000000E+1   1.000000E+1   9.000000E+1   1.100000E+1   1.100000E+1   -5.858670E-2   8.107856E-2   -8.902665E-5   -9.674329E-6   9.674329E-6   -8.902665E-5   8.955075E-5   -1.737981E+2   -8.379813E+1   
5.665866E+3   1.200117E+2   1.200117E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   -5.909904E-2   8.075184E-2   -8.913060E-5   -9.081785E-6   9.081785E-6   -8.913060E-5   8.959210E-5   -1.741820E+2   -8.418204E+1   
5.687787E+3   1.199862E+2   1.199862E+2   1.500000E+1   1.500000E+1   9.000000E+1   1.600000E+1   1.600000E+1   -5.991664E-2   8.139027E-2   -9.005189E-5   -8.894452E-6   8.894452E-6   -9.005189E-5   9.049008E-5   -1.743592E+2   -8.435917E+1   
5.709786E+3   1.199893E+2   1.199893E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   -5.809276E-2   8.046806E-2   -8.832365E-5   -9.640537E-6   9.640537E-6   -8.832365E-5   8.884823E-5   -1.737708E+2   -8.377082E+1   
5.731666E+3   1.200555E+2   1.200555E+2   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   -5.788874E-2   8.057390E-2   -8.826646E-5   -9.860625E-6   9.860625E-6   -8.826646E-5   8.881553E-5   -1.736257E+2   -8.362567E+1   
5.753516E+3   1.200535E+2   1.200535E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   -5.841920E-2   8.081688E-2   -8.875266E-5   -9.627133E-6   9.627133E-6   -8.875266E-5   8.927327E-5   -1.738092E+2   -8.380925E+1   
5.775385E+3   1.200078E+2   1.200078E+2   2.200000E+1   2.200000E+1   9.000000E+1   2.300000E+1   2.300000E+1   -5.921440E-2   7.966487E-2   -8.849399E-5   -8.285833E-6   8.285833E-6   -8.849399E-5   8.888106E-5   -1.746509E+2   -8.465090E+1   
5.797237E+3   1.201034E+2   1.201034E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   -5.977122E-2   8.104390E-2   -8.973639E-5   -8.775560E-6   8.775560E-6   -8.973639E-5   9.016447E-5   -1.744147E+2   -8.441465E+1   
5.819127E+3   1.199929E+2   1.199929E+2   2.600000E+1   2.600000E+1   9.000000E+1   2.700000E+1   2.700000E+1   -5.902327E-2   8.060734E-2   -8.898965E-5   -9.043359E-6   9.043359E-6   -8.898965E-5   8.944798E-5   -1.741974E+2   -8.419737E+1   
5.841011E+3   1.199497E+2   1.199497E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   -5.783660E-2   7.968176E-2   -8.765318E-5   -9.315936E-6   9.315936E-6   -8.765318E-5   8.814684E-5   -1.739333E+2   -8.393328E+1   
5.862992E+3   1.200409E+2   1.200409E+2   3.100000E+1   3.100000E+1   9.000000E+1   3.100000E+1   3.100000E+1   -5.913310E-2   8.097794E-2   -8.929892E-5   -9.204415E-6   9.204415E-6   -8.929892E-5   8.977204E-5   -1.741151E+2   -8.411507E+1   
5.885044E+3   1.200380E+2   1.200380E+2   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   -5.808908E-2   8.111997E-2   -8.874597E-5   -1.006946E-5   1.006946E-5   -8.874597E-5   8.931540E-5   -1.735267E+2   -8.352669E+1   
5.906939E+3   1.199986E+2   1.199986E+2   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   -5.983502E-2   8.101722E-2   -8.975847E-5   -8.710930E-6   8.710930E-6   -8.975847E-5   9.018017E-5   -1.744569E+2   -8.445689E+1   
5.928877E+3   1.199955E+2   1.199955E+2   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   -5.938712E-2   8.083221E-2   -8.936105E-5   -8.921260E-6   8.921260E-6   -8.936105E-5   8.980527E-5   -1.742988E+2   -8.429883E+1   
5.950749E+3   1.200799E+2   1.200799E+2   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   -5.888827E-2   8.141238E-2   -8.943050E-5   -9.669525E-6   9.669525E-6   -8.943050E-5   8.995174E-5   -1.738290E+2   -8.382896E+1   
5.972583E+3   1.199742E+2   1.199742E+2   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   -5.901222E-2   8.145439E-2   -8.953450E-5   -9.605304E-6   9.605304E-6   -8.953450E-5   9.004825E-5   -1.738767E+2   -8.387670E+1   
5.994466E+3   1.200329E+2   1.200329E+2   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   -5.842871E-2   8.055088E-2   -8.858529E-5   -9.446203E-6   9.446203E-6   -8.858529E-5   8.908751E-5   -1.739133E+2   -8.391332E+1   
6.016326E+3   1.200233E+2   1.200233E+2   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   -6.023171E-2   8.054629E-2   -8.969701E-5   -8.109644E-6   8.109644E-6   -8.969701E-5   9.006286E-5   -1.748338E+2   -8.483385E+1   
6.038152E+3   1.199913E+2   1.199913E+2   4.600000E+1   4.600000E+1   9.000000E+1   4.800000E+1   4.800000E+1   -5.947977E-2   8.182838E-2   -9.006713E-5   -9.504000E-6   9.504000E-6   -9.006713E-5   9.056718E-5   -1.739764E+2   -8.397637E+1   
6.060090E+3   1.200304E+2   1.200304E+2   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   -5.853454E-2   8.098346E-2   -8.893246E-5   -9.650732E-6   9.650732E-6   -8.893246E-5   8.945456E-5   -1.738066E+2   -8.380664E+1   
6.093927E+3   1.200799E+2   1.200799E+2   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   -5.944541E-2   8.326631E-2   -9.098240E-5   -1.046949E-5   1.046949E-5   -9.098240E-5   9.158279E-5   -1.734358E+2   -8.343576E+1   
6.116457E+3   1.200338E+2   1.200338E+2   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   -6.123862E-2   8.411950E-2   -9.264672E-5   -9.700965E-6   9.700965E-6   -9.264672E-5   9.315322E-5   -1.740224E+2   -8.402239E+1   
6.138592E+3   1.200368E+2   1.200368E+2   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   -6.262348E-2   8.583385E-2   -9.461944E-5   -9.797479E-6   9.797479E-6   -9.461944E-5   9.512533E-5   -1.740883E+2   -8.408831E+1   
6.160923E+3   1.200284E+2   1.200284E+2   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   -6.291124E-2   8.734327E-2   -9.578042E-5   -1.057146E-5   1.057146E-5   -9.578042E-5   9.636204E-5   -1.737017E+2   -8.370165E+1   
6.183817E+3   1.200134E+2   1.200134E+2   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   -6.377825E-2   8.845603E-2   -9.704117E-5   -1.065768E-5   1.065768E-5   -9.704117E-5   9.762466E-5   -1.737325E+2   -8.373253E+1   
6.205985E+3   1.199941E+2   1.199941E+2   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   -6.461548E-2   9.069685E-2   -9.901820E-5   -1.150342E-5   1.150342E-5   -9.901820E-5   9.968417E-5   -1.733734E+2   -8.337338E+1   
6.228125E+3   1.199830E+2   1.199830E+2   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   -6.667130E-2   9.221458E-2   -1.012777E-4   -1.097513E-5   1.097513E-5   -1.012777E-4   1.018706E-4   -1.738152E+2   -8.381518E+1   
6.250929E+3   1.200390E+2   1.200390E+2   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   -6.712782E-2   9.329947E-2   -1.022665E-4   -1.134674E-5   1.134674E-5   -1.022665E-4   1.028941E-4   -1.736688E+2   -8.366878E+1   
6.273056E+3   1.200258E+2   1.200258E+2   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   -6.918484E-2   9.541525E-2   -1.049162E-4   -1.120854E-5   1.120854E-5   -1.049162E-4   1.055133E-4   -1.739020E+2   -8.390204E+1   
6.295685E+3   1.201009E+2   1.201009E+2   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   -7.022948E-2   9.558058E-2   -1.056698E-4   -1.054398E-5   1.054398E-5   -1.056698E-4   1.061945E-4   -1.743018E+2   -8.430175E+1   
6.318593E+3   1.200009E+2   1.200009E+2   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   -7.128483E-2   9.735639E-2   -1.074788E-4   -1.092439E-5   1.092439E-5   -1.074788E-4   1.080326E-4   -1.741963E+2   -8.419626E+1   
6.341177E+3   1.200453E+2   1.200453E+2   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   -7.010829E-2   9.964356E-2   -1.082410E-4   -1.328988E-5   1.328988E-5   -1.082410E-4   1.090538E-4   -1.730002E+2   -8.300023E+1   
6.364075E+3   1.200678E+2   1.200678E+2   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   -7.182572E-2   1.016402E-1   -1.106032E-4   -1.332495E-5   1.332495E-5   -1.106032E-4   1.114030E-4   -1.731304E+2   -8.313039E+1   
6.387478E+3   1.200424E+2   1.200424E+2   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   -7.282372E-2   1.037948E-1   -1.126235E-4   -1.399541E-5   1.399541E-5   -1.126235E-4   1.134897E-4   -1.729163E+2   -8.291633E+1   
6.410153E+3   1.199390E+2   1.199390E+2   7.970000E+2   7.970000E+2   9.000000E+1   7.980000E+2   7.980000E+2   -7.352628E-2   1.047989E-1   -1.137118E-4   -1.413224E-5   1.413224E-5   -1.137118E-4   1.145866E-4   -1.729155E+2   -8.291554E+1   
6.432691E+3   1.200687E+2   1.200687E+2   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   -7.582415E-2   1.051907E-1   -1.153876E-4   -1.268879E-5   1.268879E-5   -1.153876E-4   1.160832E-4   -1.737246E+2   -8.372459E+1   
6.455952E+3   1.199686E+2   1.199686E+2   8.970000E+2   8.970000E+2   9.000000E+1   8.980000E+2   8.980000E+2   -7.620609E-2   1.062786E-1   -1.163323E-4   -1.311753E-5   1.311753E-5   -1.163323E-4   1.170695E-4   -1.735666E+2   -8.356655E+1   
6.478564E+3   1.200699E+2   1.200699E+2   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   -7.688166E-2   1.078125E-1   -1.177490E-4   -1.362072E-5   1.362072E-5   -1.177490E-4   1.185342E-4   -1.734016E+2   -8.340159E+1   
6.501149E+3   1.200579E+2   1.200579E+2   9.980000E+2   9.980000E+2   9.000000E+1   9.980000E+2   9.980000E+2   -7.837021E-2   1.108433E-1   -1.206432E-4   -1.450119E-5   1.450119E-5   -1.206432E-4   1.215116E-4   -1.731460E+2   -8.314599E+1   
6.524712E+3   1.200353E+2   1.200353E+2   1.047000E+3   1.047000E+3   9.000000E+1   1.048000E+3   1.048000E+3   -7.839016E-2   1.118472E-1   -1.213093E-4   -1.514272E-5   1.514272E-5   -1.213093E-4   1.222508E-4   -1.728847E+2   -8.288472E+1   
6.547591E+3   1.199877E+2   1.199877E+2   1.098000E+3   1.098000E+3   9.000000E+1   1.098000E+3   1.098000E+3   -8.061471E-2   1.129089E-1   -1.233762E-4   -1.419154E-5   1.419154E-5   -1.233762E-4   1.241897E-4   -1.734383E+2   -8.343830E+1   
6.570390E+3   1.200063E+2   1.200063E+2   1.148000E+3   1.148000E+3   9.000000E+1   1.148000E+3   1.148000E+3   -8.221278E-2   1.147006E-1   -1.255311E-4   -1.418091E-5   1.418091E-5   -1.255311E-4   1.263295E-4   -1.735548E+2   -8.355477E+1   
6.593928E+3   1.200460E+2   1.200460E+2   1.197000E+3   1.197000E+3   9.000000E+1   1.198000E+3   1.198000E+3   -8.246989E-2   1.154372E-1   -1.261698E-4   -1.447232E-5   1.447232E-5   -1.261698E-4   1.269971E-4   -1.734565E+2   -8.345648E+1   
6.616770E+3   1.200015E+2   1.200015E+2   1.248000E+3   1.248000E+3   9.000000E+1   1.248000E+3   1.248000E+3   -8.313652E-2   1.171672E-1   -1.277087E-4   -1.511028E-5   1.511028E-5   -1.277087E-4   1.285995E-4   -1.732522E+2   -8.325223E+1   
6.639583E+3   1.200255E+2   1.200255E+2   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   -8.140132E-2   1.182380E-1   -1.273332E-4   -1.709369E-5   1.709369E-5   -1.273332E-4   1.284755E-4   -1.723541E+2   -8.235411E+1   
6.663164E+3   1.200784E+2   1.200784E+2   1.348000E+3   1.348000E+3   9.000000E+1   1.348000E+3   1.348000E+3   -8.344979E-2   1.191767E-1   -1.292111E-4   -1.619233E-5   1.619233E-5   -1.292111E-4   1.302217E-4   -1.728571E+2   -8.285711E+1   
6.685744E+3   1.200515E+2   1.200515E+2   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   -8.574522E-2   1.202505E-1   -1.313296E-4   -1.519656E-5   1.519656E-5   -1.313296E-4   1.322059E-4   -1.733995E+2   -8.339948E+1   
6.708277E+3   1.199872E+2   1.199872E+2   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   -8.685027E-2   1.229432E-1   -1.337665E-4   -1.613966E-5   1.613966E-5   -1.337665E-4   1.347367E-4   -1.731202E+2   -8.312021E+1   
6.731272E+3   1.199816E+2   1.199816E+2   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   -8.761172E-2   1.234991E-1   -1.345993E-4   -1.593990E-5   1.593990E-5   -1.345993E-4   1.355399E-4   -1.732462E+2   -8.324622E+1   
6.753860E+3   1.200020E+2   1.200020E+2   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   -8.717546E-2   1.262011E-1   -1.360894E-4   -1.802901E-5   1.802901E-5   -1.360894E-4   1.372784E-4   -1.724534E+2   -8.245344E+1   
6.776395E+3   1.200860E+2   1.200860E+2   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   -8.955897E-2   1.266410E-1   -1.378495E-4   -1.655371E-5   1.655371E-5   -1.378495E-4   1.388399E-4   -1.731524E+2   -8.315240E+1   
6.799681E+3   1.200671E+2   1.200671E+2   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   -9.034771E-2   1.281523E-1   -1.393214E-4   -1.695836E-5   1.695836E-5   -1.393214E-4   1.403497E-4   -1.730600E+2   -8.306003E+1   
6.822229E+3   1.199830E+2   1.199830E+2   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   -9.116596E-2   1.298034E-1   -1.409026E-4   -1.743263E-5   1.743263E-5   -1.409026E-4   1.419769E-4   -1.729471E+2   -8.294714E+1   
6.844809E+3   1.200394E+2   1.200394E+2   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   -9.273773E-2   1.316552E-1   -1.430805E-4   -1.748076E-5   1.748076E-5   -1.430805E-4   1.441443E-4   -1.730344E+2   -8.303445E+1   
6.867585E+3   1.199720E+2   1.199720E+2   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   -9.305093E-2   1.324737E-1   -1.438072E-4   -1.778424E-5   1.778424E-5   -1.438072E-4   1.449027E-4   -1.729502E+2   -8.295018E+1   
6.890136E+3   1.199516E+2   1.199516E+2   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   -9.252942E-2   1.338884E-1   -1.444061E-4   -1.909480E-5   1.909480E-5   -1.444061E-4   1.456631E-4   -1.724675E+2   -8.246748E+1   
6.912719E+3   1.200515E+2   1.200515E+2   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   -9.493754E-2   1.376935E-1   -1.483732E-4   -1.980137E-5   1.980137E-5   -1.483732E-4   1.496886E-4   -1.723984E+2   -8.239842E+1   
6.935548E+3   1.200576E+2   1.200576E+2   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   -9.708272E-2   1.381071E-1   -1.499687E-4   -1.848511E-5   1.848511E-5   -1.499687E-4   1.511037E-4   -1.729732E+2   -8.297318E+1   
6.958087E+3   1.199894E+2   1.199894E+2   1.999000E+3   1.999000E+3   9.000000E+1   2.000000E+3   2.000000E+3   -9.766901E-2   1.401641E-1   -1.516709E-4   -1.939630E-5   1.939630E-5   -1.516709E-4   1.529062E-4   -1.727123E+2   -8.271234E+1   
6.996041E+3   1.199788E+2   1.199788E+2   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   -1.110777E-1   1.567269E-1   -1.707480E-4   -2.030711E-5   2.030711E-5   -1.707480E-4   1.719514E-4   -1.732177E+2   -8.321766E+1   
7.022471E+3   1.199992E+2   1.199992E+2   2.998000E+3   2.998000E+3   9.000000E+1   2.998000E+3   2.998000E+3   -1.221376E-1   1.753250E-1   -1.896985E-4   -2.428576E-5   2.428576E-5   -1.896985E-4   1.912467E-4   -1.727045E+2   -8.270451E+1   
7.048372E+3   1.200824E+2   1.200824E+2   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -1.357687E-1   1.930951E-1   -2.096994E-4   -2.582140E-5   2.582140E-5   -2.096994E-4   2.112832E-4   -1.729802E+2   -8.298020E+1   
7.074177E+3   1.200232E+2   1.200232E+2   3.998000E+3   3.998000E+3   9.000000E+1   4.000000E+3   4.000000E+3   -1.448215E-1   2.077789E-1   -2.248596E-4   -2.872545E-5   2.872545E-5   -2.248596E-4   2.266870E-4   -1.727200E+2   -8.271999E+1   
7.100684E+3   1.199738E+2   1.199738E+2   4.498000E+3   4.498000E+3   9.000000E+1   4.499000E+3   4.499000E+3   -1.463058E-1   2.144034E-1   -2.300918E-4   -3.195858E-5   3.195858E-5   -2.300918E-4   2.323006E-4   -1.720925E+2   -8.209250E+1   
7.126905E+3   1.200305E+2   1.200305E+2   4.998000E+3   4.998000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -1.432627E-1   2.120371E-1   -2.266692E-4   -3.266233E-5   3.266233E-5   -2.266692E-4   2.290104E-4   -1.718003E+2   -8.180030E+1   
7.152537E+3   1.200693E+2   1.200693E+2   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -1.288054E-1   1.965417E-1   -2.076390E-4   -3.322489E-5   3.322489E-5   -2.076390E-4   2.102804E-4   -1.709090E+2   -8.090901E+1   
7.178984E+3   1.199957E+2   1.199957E+2   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -1.118696E-1   1.795983E-1   -1.861335E-4   -3.467410E-5   3.467410E-5   -1.861335E-4   1.893356E-4   -1.694475E+2   -7.944754E+1   
7.204927E+3   1.200709E+2   1.200709E+2   6.497000E+3   6.497000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -1.019295E-1   1.690235E-1   -1.731008E-4   -3.511256E-5   3.511256E-5   -1.731008E-4   1.766261E-4   -1.685334E+2   -7.853344E+1   
7.231151E+3   1.199719E+2   1.199719E+2   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -9.466016E-2   1.628352E-1   -1.645762E-4   -3.644345E-5   3.644345E-5   -1.645762E-4   1.685629E-4   -1.675140E+2   -7.751401E+1   
7.256826E+3   1.200290E+2   1.200290E+2   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -9.851238E-2   1.691898E-1   -1.710965E-4   -3.774867E-5   3.774867E-5   -1.710965E-4   1.752112E-4   -1.675583E+2   -7.755826E+1   
7.282260E+3   1.200618E+2   1.200618E+2   7.999000E+3   7.999000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -1.011382E-1   1.761340E-1   -1.772426E-4   -4.034645E-5   4.034645E-5   -1.772426E-4   1.817767E-4   -1.671760E+2   -7.717605E+1   
7.308672E+3   1.200518E+2   1.200518E+2   8.498000E+3   8.498000E+3   9.000000E+1   8.499000E+3   8.499000E+3   -1.136345E-1   1.920709E-1   -1.953480E-4   -4.152292E-5   4.152292E-5   -1.953480E-4   1.997122E-4   -1.679999E+2   -7.799988E+1   
7.335076E+3   1.200025E+2   1.200025E+2   8.998000E+3   8.998000E+3   9.000000E+1   8.999000E+3   8.999000E+3   -1.249840E-1   2.091867E-1   -2.135121E-4   -4.431832E-5   4.431832E-5   -2.135121E-4   2.180631E-4   -1.682737E+2   -7.827373E+1   
7.361469E+3   1.200523E+2   1.200523E+2   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -1.338160E-1   2.252136E-1   -2.294105E-4   -4.826383E-5   4.826383E-5   -2.294105E-4   2.344324E-4   -1.681193E+2   -7.811926E+1   
7.387377E+3   1.200825E+2   1.200825E+2   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -1.453210E-1   2.420737E-1   -2.475042E-4   -5.077700E-5   5.077700E-5   -2.475042E-4   2.526592E-4   -1.684063E+2   -7.840629E+1   
@@END Data.
@Time at end of measurement: 15:12:44
@NO Instrument  Changes.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -9499.000      -9999.000      250.000        Coercive Field: Field at which M//H changes sign
Ms  emu                                 3.179E-4       -3.114E-4      3.146E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -8.870E-5      1.346E-4       1.116E-4       Remanent Magnetization: M at H=0        
S                                       0.279          0.432          0.356          Squareness: Mr/Ms                       
S*                                      1.636          1.166          1.401          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
