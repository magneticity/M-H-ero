@Filename: c:\vsm-lv\Will\data\AJA901_700sNiFe_on_CoPd8\AJA901_700sNiFe_on_CoPd8_outOfPlane_loop.VHD
@Measurement Controlfilename: c:\vsm-lv\Will\Recipes\full20000GaussHys_outOfPlane.VHC
@Signal Manipulation filename: c:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA901_700sNiFe_on_CoPd8
@Date: 08 March 2019    (2019-08-03)
@Time: 11:41:03
@Test ID: AJA901_700sNiFe_on_CoPd8_outOfPlaneLoop
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 89.9995 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Applied Field to 19997.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Auto Range Signal to 13.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 4
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 5.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 20000.0000 [Oe] To: 5000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 5000.0000 [Oe] To:  0.0000 [Oe] Min Stepsize/Sweeprate = 200.0000 [Oe] Max Stepsize/Sweeprate = 200.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From:  0.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 200.0000 [Oe] Max Stepsize/Sweeprate = 200.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -20000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 3 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 50 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 25.915
@Y Coils Correction Factor: 0.996
@Sample Shape Correction Factor: 0.896
@Coil Angle Alpha: 41.920
@Coil Angle Beta: -48.000
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
15000.000000   1.000000
15249.000000   1.000524
15499.000000   1.000702
15750.000000   1.001233
16000.000000   1.001406
16250.000000   1.001585
16499.000000   1.001758
16749.000000   1.001937
16999.000000   1.002110
17249.000000   1.001937
17499.000000   1.002289
17749.000000   1.002289
17999.000000   1.002289
18249.000000   1.002462
18499.000000   1.002462
18748.000000   1.002462
18999.000000   1.002462
19249.000000   1.002462
19499.000000   1.002642
19749.000000   1.002642
19999.000000   1.002462
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = No
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 03 December 2018  15:19:40
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 4
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 11:41:03
@@Data
New Section: Section 0: 
3.295900E+1   2.148089E+1   2.148089E+1   1.999700E+4   1.999700E+4   8.999955E+1   1.999700E+4   1.999700E+4   -4.485590E-1   5.977000E-1   -6.660931E-4   -6.447056E-5   6.446533E-5   -6.660936E-4   6.692058E-4   -1.744716E+2   -8.447206E+1   
6.136300E+1   2.148419E+1   2.148419E+1   1.949700E+4   1.949700E+4   8.999955E+1   1.949700E+4   1.949700E+4   -4.186363E-1   5.640690E-1   -6.259153E-4   -6.432785E-5   6.432293E-5   -6.259158E-4   6.292122E-4   -1.741321E+2   -8.413253E+1   
8.921500E+1   2.150341E+1   2.150341E+1   1.899600E+4   1.899600E+4   8.999955E+1   1.899600E+4   1.899600E+4   -3.870915E-1   5.289985E-1   -5.835863E-4   -6.443301E-5   6.442842E-5   -5.835868E-4   5.871325E-4   -1.736996E+2   -8.370002E+1   
1.166140E+2   2.149911E+1   2.149911E+1   1.849600E+4   1.849600E+4   8.999955E+1   1.849700E+4   1.849700E+4   -3.583636E-1   4.968643E-1   -5.450089E-4   -6.439848E-5   6.439420E-5   -5.450094E-4   5.488004E-4   -1.732612E+2   -8.326160E+1   
1.433590E+2   2.148651E+1   2.148651E+1   1.799700E+4   1.799700E+4   8.999955E+1   1.799700E+4   1.799700E+4   -3.214957E-1   4.589892E-1   -4.976497E-4   -6.659581E-5   6.659190E-5   -4.976502E-4   5.020859E-4   -1.723779E+2   -8.237837E+1   
1.698970E+2   2.146520E+1   2.146520E+1   1.749700E+4   1.749700E+4   8.999955E+1   1.749700E+4   1.749700E+4   -2.937482E-1   4.293901E-1   -4.613494E-4   -6.752083E-5   6.751721E-5   -4.613500E-4   4.662643E-4   -1.716736E+2   -8.167404E+1   
1.967970E+2   2.146639E+1   2.146639E+1   1.699600E+4   1.699600E+4   8.999955E+1   1.699600E+4   1.699600E+4   -2.660136E-1   3.986943E-1   -4.242543E-4   -6.770566E-5   6.770233E-5   -4.242548E-4   4.296228E-4   -1.709328E+2   -8.093322E+1   
2.229950E+2   2.144390E+1   2.144390E+1   1.649700E+4   1.649700E+4   8.999955E+1   1.649700E+4   1.649700E+4   -2.340744E-1   3.659884E-1   -3.832511E-4   -6.967966E-5   6.967665E-5   -3.832517E-4   3.895339E-4   -1.696955E+2   -7.969595E+1   
2.491880E+2   2.143200E+1   2.143200E+1   1.599700E+4   1.599700E+4   8.999955E+1   1.599800E+4   1.599800E+4   -1.963907E-1   3.286010E-1   -3.357278E-4   -7.280892E-5   7.280629E-5   -3.357284E-4   3.435321E-4   -1.677638E+2   -7.776426E+1   
2.746360E+2   2.143560E+1   2.143560E+1   1.549600E+4   1.549600E+4   8.999955E+1   1.549700E+4   1.549700E+4   -1.721891E-1   3.005253E-1   -3.023836E-4   -7.211063E-5   7.210825E-5   -3.023842E-4   3.108630E-4   -1.665870E+2   -7.658742E+1   
3.002610E+2   2.140591E+1   2.140591E+1   1.499700E+4   1.499700E+4   8.999955E+1   1.499700E+4   1.499700E+4   -1.405073E-1   2.715757E-1   -2.640322E-4   -7.639581E-5   7.639373E-5   -2.640328E-4   2.748624E-4   -1.638626E+2   -7.386303E+1   
3.256490E+2   2.136639E+1   2.136639E+1   1.449700E+4   1.449700E+4   8.999955E+1   1.449700E+4   1.449700E+4   -1.080094E-1   2.386852E-1   -2.227927E-4   -7.866259E-5   7.866084E-5   -2.227934E-4   2.362719E-4   -1.605531E+2   -7.055359E+1   
3.508470E+2   2.137289E+1   2.137289E+1   1.399700E+4   1.399700E+4   8.999955E+1   1.399700E+4   1.399700E+4   -7.343240E-2   2.063913E-1   -1.807047E-4   -8.287390E-5   8.287248E-5   -1.807054E-4   1.988021E-4   -1.553631E+2   -6.536355E+1   
3.763490E+2   2.139700E+1   2.139700E+1   1.349700E+4   1.349700E+4   8.999955E+1   1.349700E+4   1.349700E+4   -4.111522E-2   1.754921E-1   -1.408929E-4   -8.633292E-5   8.633181E-5   -1.408936E-4   1.652398E-4   -1.485019E+2   -5.850233E+1   
4.015340E+2   2.138229E+1   2.138229E+1   1.299600E+4   1.299600E+4   8.999955E+1   1.299600E+4   1.299600E+4   -1.170648E-2   1.482093E-1   -1.052178E-4   -9.003739E-5   9.003656E-5   -1.052185E-4   1.384829E-4   -1.394456E+2   -4.944606E+1   
4.270260E+2   2.143649E+1   2.143649E+1   1.249700E+4   1.249700E+4   8.999955E+1   1.249700E+4   1.249700E+4   2.152269E-2   1.211048E-1   -6.737501E-5   -9.670333E-5   9.670280E-5   -6.737577E-5   1.178598E-4   -1.248656E+2   -3.486610E+1   
4.519670E+2   2.145849E+1   2.145849E+1   1.199700E+4   1.199700E+4   8.999955E+1   1.199700E+4   1.199700E+4   5.803813E-2   9.292962E-2   -2.685653E-5   -1.051012E-4   1.051010E-4   -2.685736E-5   1.084782E-4   -1.043341E+2   -1.433453E+1   
4.774520E+2   2.147000E+1   2.147000E+1   1.149700E+4   1.149700E+4   8.999955E+1   1.149700E+4   1.149700E+4   9.369749E-2   7.023115E-2   9.520521E-6   -1.165110E-4   1.165110E-4   9.519606E-6   1.168993E-4   -8.532854E+1   4.671011E+0   
5.026330E+2   2.146801E+1   2.146801E+1   1.099600E+4   1.099600E+4   8.999955E+1   1.099600E+4   1.099600E+4   1.309106E-1   4.739678E-2   4.691728E-5   -1.289864E-4   1.289867E-4   4.691627E-5   1.372542E-4   -7.001173E+1   1.998782E+1   
5.276180E+2   2.146938E+1   2.146938E+1   1.049700E+4   1.049700E+4   8.999955E+1   1.049700E+4   1.049700E+4   1.697409E-1   2.989791E-2   8.174591E-5   -1.462199E-4   1.462205E-4   8.174476E-5   1.675191E-4   -6.079212E+1   2.920743E+1   
5.526640E+2   2.147369E+1   2.147369E+1   9.997000E+3   9.997000E+3   8.999955E+1   9.997000E+3   9.997000E+3   2.102600E-1   1.900878E-2   1.132050E-4   -1.691140E-4   1.691149E-4   1.132036E-4   2.035065E-4   -5.620163E+1   3.379792E+1   
5.778080E+2   2.148870E+1   2.148870E+1   9.497000E+3   9.497000E+3   8.999955E+1   9.497000E+3   9.497000E+3   2.522130E-1   1.310953E-2   1.422152E-4   -1.963996E-4   1.964007E-4   1.422137E-4   2.424829E-4   -5.409126E+1   3.590829E+1   
6.029080E+2   2.148620E+1   2.148620E+1   8.996000E+3   8.996000E+3   8.999955E+1   8.997000E+3   8.997000E+3   2.979606E-1   1.130680E-2   1.707813E-4   -2.292380E-4   2.292394E-4   1.707795E-4   2.858607E-4   -5.331406E+1   3.668549E+1   
6.279990E+2   2.151251E+1   2.151251E+1   8.496000E+3   8.496000E+3   8.999955E+1   8.497000E+3   8.497000E+3   3.397128E-1   1.706639E-2   1.919455E-4   -2.641422E-4   2.641437E-4   1.919435E-4   3.265183E-4   -5.399504E+1   3.600451E+1   
6.530770E+2   2.151660E+1   2.151660E+1   7.997000E+3   7.997000E+3   8.999955E+1   7.998000E+3   7.998000E+3   3.822971E-1   2.760926E-2   2.104379E-4   -3.028525E-4   3.028542E-4   2.104355E-4   3.687869E-4   -5.520639E+1   3.479316E+1   
6.784220E+2   2.152770E+1   2.152770E+1   7.497000E+3   7.497000E+3   8.999955E+1   7.497000E+3   7.497000E+3   4.222144E-1   3.731603E-2   2.278886E-4   -3.390213E-4   3.390231E-4   2.278859E-4   4.084956E-4   -5.609118E+1   3.390837E+1   
7.037410E+2   2.153939E+1   2.153939E+1   6.996000E+3   6.996000E+3   8.999955E+1   6.996000E+3   6.996000E+3   4.568181E-1   5.287517E-2   2.382819E-4   -3.751357E-4   3.751375E-4   2.382790E-4   4.444154E-4   -5.757675E+1   3.242280E+1   
7.288430E+2   2.153439E+1   2.153439E+1   6.496000E+3   6.496000E+3   8.999955E+1   6.497000E+3   6.497000E+3   4.876442E-1   6.611790E-2   2.479501E-4   -4.068958E-4   4.068978E-4   2.479469E-4   4.764908E-4   -5.864313E+1   3.135642E+1   
7.536350E+2   2.154391E+1   2.154391E+1   5.996000E+3   5.996000E+3   8.999955E+1   5.997000E+3   5.997000E+3   5.193683E-1   7.823815E-2   2.588993E-4   -4.385763E-4   4.385783E-4   2.588959E-4   5.092916E-4   -5.944590E+1   3.055365E+1   
7.790170E+2   2.154461E+1   2.154461E+1   5.496000E+3   5.496000E+3   8.999955E+1   5.497000E+3   5.497000E+3   5.482305E-1   9.156839E-2   2.673344E-4   -4.689334E-4   4.689355E-4   2.673307E-4   5.397835E-4   -6.031295E+1   2.968660E+1   
8.041220E+2   2.157501E+1   2.157501E+1   4.996000E+3   4.996000E+3   8.999955E+1   4.996000E+3   4.996000E+3   5.700832E-1   1.061604E-1   2.707395E-4   -4.949158E-4   4.949179E-4   2.707357E-4   5.641290E-4   -6.131950E+1   2.868005E+1   
8.391610E+2   2.159191E+1   2.159191E+1   4.796000E+3   4.796000E+3   8.999955E+1   4.797000E+3   4.797000E+3   5.806549E-1   1.090251E-1   2.751664E-4   -5.046905E-4   5.046927E-4   2.751625E-4   5.748296E-4   -6.139998E+1   2.859957E+1   
8.628870E+2   2.159249E+1   2.159249E+1   4.596000E+3   4.596000E+3   8.999955E+1   4.596000E+3   4.596000E+3   5.900277E-1   1.137594E-1   2.776370E-4   -5.148189E-4   5.148211E-4   2.776330E-4   5.849110E-4   -6.166243E+1   2.833712E+1   
8.866170E+2   2.159731E+1   2.159731E+1   4.397000E+3   4.397000E+3   8.999955E+1   4.397000E+3   4.397000E+3   5.987305E-1   1.192776E-1   2.791873E-4   -5.249711E-4   5.249733E-4   2.791831E-4   5.945924E-4   -6.199530E+1   2.800425E+1   
9.100670E+2   2.160571E+1   2.160571E+1   4.197000E+3   4.197000E+3   8.999955E+1   4.197000E+3   4.197000E+3   6.072870E-1   1.245229E-1   2.808309E-4   -5.348326E-4   5.348348E-4   2.808267E-4   6.040794E-4   -6.229685E+1   2.770270E+1   
9.337380E+2   2.159930E+1   2.159930E+1   3.997000E+3   3.997000E+3   8.999955E+1   3.998000E+3   3.998000E+3   6.154506E-1   1.288524E-1   2.828462E-4   -5.437915E-4   5.437937E-4   2.828419E-4   6.129528E-4   -6.251938E+1   2.748017E+1   
9.574070E+2   2.161050E+1   2.161050E+1   3.797000E+3   3.797000E+3   8.999955E+1   3.798000E+3   3.798000E+3   6.251581E-1   1.321605E-1   2.864621E-4   -5.532187E-4   5.532209E-4   2.864578E-4   6.229859E-4   -6.262443E+1   2.737512E+1   
9.808850E+2   2.162328E+1   2.162328E+1   3.597000E+3   3.597000E+3   8.999955E+1   3.597000E+3   3.597000E+3   6.310798E-1   1.385656E-1   2.857608E-4   -5.618924E-4   5.618947E-4   2.857563E-4   6.303827E-4   -6.304355E+1   2.695600E+1   
1.004581E+3   2.162231E+1   2.162231E+1   3.397000E+3   3.397000E+3   8.999955E+1   3.397000E+3   3.397000E+3   6.379399E-1   1.420281E-1   2.875707E-4   -5.693038E-4   5.693061E-4   2.875662E-4   6.378117E-4   -6.320043E+1   2.679912E+1   
1.028011E+3   2.163311E+1   2.163311E+1   3.197000E+3   3.197000E+3   8.999955E+1   3.197000E+3   3.197000E+3   6.468182E-1   1.466003E-1   2.898529E-4   -5.789562E-4   5.789585E-4   2.898484E-4   6.474604E-4   -6.340528E+1   2.659427E+1   
1.051649E+3   2.163149E+1   2.163149E+1   2.996000E+3   2.996000E+3   8.999955E+1   2.997000E+3   2.997000E+3   6.533360E-1   1.513294E-1   2.906187E-4   -5.869569E-4   5.869591E-4   2.906141E-4   6.549638E-4   -6.365870E+1   2.634085E+1   
1.075392E+3   2.161950E+1   2.161950E+1   2.797000E+3   2.797000E+3   8.999955E+1   2.797000E+3   2.797000E+3   6.604825E-1   1.554247E-1   2.921808E-4   -5.950029E-4   5.950052E-4   2.921761E-4   6.628711E-4   -6.384630E+1   2.615325E+1   
1.099001E+3   2.167321E+1   2.167321E+1   2.596000E+3   2.596000E+3   8.999955E+1   2.597000E+3   2.597000E+3   6.671089E-1   1.610253E-1   2.924341E-4   -6.036650E-4   6.036673E-4   2.924294E-4   6.707676E-4   -6.415301E+1   2.584654E+1   
1.122617E+3   2.166830E+1   2.166830E+1   2.397000E+3   2.397000E+3   8.999955E+1   2.397000E+3   2.397000E+3   6.732143E-1   1.635597E-1   2.944076E-4   -6.098965E-4   6.098989E-4   2.944028E-4   6.772367E-4   -6.423260E+1   2.576695E+1   
1.146269E+3   2.167831E+1   2.167831E+1   2.197000E+3   2.197000E+3   8.999955E+1   2.198000E+3   2.198000E+3   6.804185E-1   1.691172E-1   2.950352E-4   -6.189598E-4   6.189621E-4   2.950303E-4   6.856800E-4   -6.451459E+1   2.548496E+1   
1.169913E+3   2.169271E+1   2.169271E+1   1.997000E+3   1.997000E+3   8.999955E+1   1.998000E+3   1.998000E+3   6.863159E-1   1.730103E-1   2.959838E-4   -6.259418E-4   6.259441E-4   2.959789E-4   6.923940E-4   -6.469233E+1   2.530722E+1   
1.193317E+3   2.167971E+1   2.167971E+1   1.797000E+3   1.797000E+3   8.999955E+1   1.797000E+3   1.797000E+3   6.939543E-1   1.780278E-1   2.972290E-4   -6.349683E-4   6.349706E-4   2.972240E-4   7.010919E-4   -6.491568E+1   2.508387E+1   
1.216789E+3   2.168401E+1   2.168401E+1   1.597000E+3   1.597000E+3   8.999955E+1   1.597000E+3   1.597000E+3   7.003335E-1   1.820664E-1   2.983695E-4   -6.424057E-4   6.424080E-4   2.983645E-4   7.083145E-4   -6.508718E+1   2.491237E+1   
1.240255E+3   2.168441E+1   2.168441E+1   1.397000E+3   1.397000E+3   8.999955E+1   1.397000E+3   1.397000E+3   7.055165E-1   1.886305E-1   2.971208E-4   -6.506357E-4   6.506380E-4   2.971157E-4   7.152675E-4   -6.545561E+1   2.454394E+1   
1.263919E+3   2.167611E+1   2.167611E+1   1.197000E+3   1.197000E+3   8.999955E+1   1.197000E+3   1.197000E+3   7.145131E-1   1.945014E-1   2.986132E-4   -6.612415E-4   6.612438E-4   2.986080E-4   7.255413E-4   -6.569632E+1   2.430323E+1   
1.287447E+3   2.166729E+1   2.166729E+1   9.960000E+2   9.960000E+2   8.999955E+1   9.960000E+2   9.960000E+2   7.208276E-1   2.013062E-1   2.978818E-4   -6.704738E-4   6.704761E-4   2.978766E-4   7.336680E-4   -6.604511E+1   2.395444E+1   
1.310625E+3   2.166549E+1   2.166549E+1   7.960000E+2   7.960000E+2   8.999955E+1   7.970000E+2   7.970000E+2   7.291776E-1   2.101248E-1   2.970339E-4   -6.825624E-4   6.825647E-4   2.970286E-4   7.443928E-4   -6.648254E+1   2.351701E+1   
1.333614E+3   2.167101E+1   2.167101E+1   5.960000E+2   5.960000E+2   8.999955E+1   5.970000E+2   5.970000E+2   7.384886E-1   2.203536E-1   2.958266E-4   -6.963056E-4   6.963079E-4   2.958211E-4   7.565414E-4   -6.698171E+1   2.301784E+1   
1.356741E+3   2.167950E+1   2.167950E+1   3.970000E+2   3.970000E+2   8.999955E+1   3.970000E+2   3.970000E+2   7.513337E-1   2.345996E-1   2.940716E-4   -7.153551E-4   7.153574E-4   2.940660E-4   7.734410E-4   -6.765318E+1   2.234637E+1   
1.379542E+3   2.167571E+1   2.167571E+1   1.970000E+2   1.970000E+2   8.999955E+1   1.970000E+2   1.970000E+2   7.641456E-1   2.490175E-1   2.921828E-4   -7.344943E-4   7.344966E-4   2.921771E-4   7.904763E-4   -6.830727E+1   2.169228E+1   
1.401522E+3   2.167080E+1   2.167080E+1   -1.000000E+0   -1.000000E+0   8.999955E+1   0.000000E+0   0.000000E+0   7.509640E-1   2.478783E-1   2.850510E-4   -7.239273E-4   7.239295E-4   2.850453E-4   7.780262E-4   -6.850764E+1   2.149191E+1   
1.435821E+3   2.165890E+1   2.165890E+1   -2.010000E+2   -2.010000E+2   8.999955E+1   -2.010000E+2   -2.010000E+2   3.724378E-1   -4.126387E-2   2.501790E-4   -2.496282E-4   2.496302E-4   2.501771E-4   3.534173E-4   -4.493685E+1   4.506270E+1   
1.458511E+3   2.165789E+1   2.165789E+1   -4.010000E+2   -4.010000E+2   8.999955E+1   -4.010000E+2   -4.010000E+2   -1.470540E-1   -2.235419E-1   6.014980E-5   2.583591E-4   -2.583586E-4   6.015182E-5   2.652685E-4   7.689416E+1   1.668937E+2   
1.481681E+3   2.165359E+1   2.165359E+1   -6.010000E+2   -6.010000E+2   8.999955E+1   -6.010000E+2   -6.010000E+2   -3.710630E-1   -1.674439E-1   -1.110523E-4   3.876616E-4   -3.876625E-4   -1.110493E-4   4.032544E-4   1.059853E+2   1.959848E+2   
1.504375E+3   2.165151E+1   2.165151E+1   -8.010000E+2   -8.010000E+2   8.999955E+1   -8.010000E+2   -8.010000E+2   -5.300424E-1   -1.845211E-1   -1.948554E-4   5.173321E-4   -5.173336E-4   -1.948513E-4   5.528120E-4   1.106391E+2   2.006387E+2   
1.527051E+3   2.164550E+1   2.164550E+1   -1.001000E+3   -1.001000E+3   8.999955E+1   -1.001000E+3   -1.001000E+3   -6.406398E-1   -1.893294E-1   -2.578410E-4   6.028283E-4   -6.028303E-4   -2.578363E-4   6.556554E-4   1.131573E+2   2.031569E+2   
1.550386E+3   2.164071E+1   2.164071E+1   -1.202000E+3   -1.202000E+3   8.999955E+1   -1.201000E+3   -1.201000E+3   -6.986851E-1   -1.722683E-1   -3.038762E-4   6.346510E-4   -6.346533E-4   -3.038712E-4   7.036495E-4   1.155855E+2   2.055850E+2   
1.573225E+3   2.162802E+1   2.162802E+1   -1.401000E+3   -1.401000E+3   8.999955E+1   -1.401000E+3   -1.401000E+3   -7.087054E-1   -1.664199E-1   -3.137471E-4   6.382102E-4   -6.382127E-4   -3.137421E-4   7.111606E-4   1.161789E+2   2.061785E+2   
1.596025E+3   2.162371E+1   2.162371E+1   -1.601000E+3   -1.601000E+3   8.999955E+1   -1.600000E+3   -1.600000E+3   -7.067966E-1   -1.619404E-1   -3.155733E-4   6.338053E-4   -6.338078E-4   -3.155684E-4   7.080224E-4   1.164688E+2   2.064684E+2   
1.619776E+3   2.162328E+1   2.162328E+1   -1.801000E+3   -1.801000E+3   8.999955E+1   -1.800000E+3   -1.800000E+3   -7.061278E-1   -1.598977E-1   -3.165269E-4   6.319467E-4   -6.319492E-4   -3.165220E-4   7.067856E-4   1.166052E+2   2.066047E+2   
1.643007E+3   2.162829E+1   2.162829E+1   -2.001000E+3   -2.001000E+3   8.999955E+1   -2.000000E+3   -2.000000E+3   -7.016175E-1   -1.562272E-1   -3.162606E-4   6.261451E-4   -6.261476E-4   -3.162557E-4   7.014830E-4   1.167980E+2   2.067975E+2   
1.679009E+3   2.160610E+1   2.160610E+1   -2.501000E+3   -2.501000E+3   8.999955E+1   -2.501000E+3   -2.501000E+3   -6.873752E-1   -1.463222E-1   -3.143030E-4   6.089484E-4   -6.089509E-4   -3.142982E-4   6.852770E-4   1.173001E+2   2.072996E+2   
1.703669E+3   2.160781E+1   2.160781E+1   -3.001000E+3   -3.001000E+3   8.999955E+1   -3.001000E+3   -3.001000E+3   -6.747331E-1   -1.364025E-1   -3.133125E-4   5.929324E-4   -5.929349E-4   -3.133079E-4   6.706218E-4   1.178525E+2   2.078521E+2   
1.727867E+3   2.161120E+1   2.161120E+1   -3.501000E+3   -3.501000E+3   8.999955E+1   -3.501000E+3   -3.501000E+3   -6.565863E-1   -1.248730E-1   -3.100952E-4   5.717481E-4   -5.717506E-4   -3.100908E-4   6.504268E-4   1.184738E+2   2.084733E+2   
1.752599E+3   2.160900E+1   2.160900E+1   -4.000000E+3   -4.000000E+3   8.999955E+1   -4.000000E+3   -4.000000E+3   -6.374629E-1   -1.133925E-1   -3.062613E-4   5.498697E-4   -5.498722E-4   -3.062569E-4   6.294066E-4   1.191165E+2   2.091161E+2   
1.777291E+3   2.159219E+1   2.159219E+1   -4.501000E+3   -4.501000E+3   8.999955E+1   -4.501000E+3   -4.501000E+3   -6.142038E-1   -1.011911E-1   -3.004305E-4   5.244338E-4   -5.244361E-4   -3.004264E-4   6.043917E-4   1.198069E+2   2.098065E+2   
1.801638E+3   2.159081E+1   2.159081E+1   -5.001000E+3   -5.001000E+3   8.999955E+1   -5.001000E+3   -5.001000E+3   -5.928275E-1   -8.836196E-2   -2.961422E-4   4.999806E-4   -4.999829E-4   -2.961383E-4   5.811031E-4   1.206386E+2   2.106381E+2   
1.825852E+3   2.157711E+1   2.157711E+1   -5.501000E+3   -5.501000E+3   8.999955E+1   -5.501000E+3   -5.501000E+3   -5.701277E-1   -7.546293E-2   -2.911084E-4   4.744959E-4   -4.744982E-4   -2.911047E-4   5.566781E-4   1.215296E+2   2.115291E+2   
1.850604E+3   2.157400E+1   2.157400E+1   -6.001000E+3   -6.001000E+3   8.999955E+1   -6.001000E+3   -6.001000E+3   -5.404482E-1   -6.382088E-2   -2.810656E-4   4.446554E-4   -4.446576E-4   -2.810621E-4   5.260383E-4   1.222969E+2   2.122964E+2   
1.874813E+3   2.155499E+1   2.155499E+1   -6.502000E+3   -6.502000E+3   8.999955E+1   -6.501000E+3   -6.501000E+3   -5.118769E-1   -4.885326E-2   -2.738895E-4   4.134237E-4   -4.134259E-4   -2.738863E-4   4.959180E-4   1.235241E+2   2.135237E+2   
1.898610E+3   2.156140E+1   2.156140E+1   -7.002000E+3   -7.002000E+3   8.999955E+1   -7.002000E+3   -7.002000E+3   -4.780211E-1   -3.734950E-2   -2.612563E-4   3.805679E-4   -3.805699E-4   -2.612533E-4   4.616133E-4   1.244692E+2   2.144688E+2   
1.922801E+3   2.154781E+1   2.154781E+1   -7.501000E+3   -7.501000E+3   8.999955E+1   -7.501000E+3   -7.501000E+3   -4.401337E-1   -2.442277E-2   -2.471539E-4   3.437642E-4   -3.437661E-4   -2.471512E-4   4.233897E-4   1.257148E+2   2.157143E+2   
1.947073E+3   2.154049E+1   2.154049E+1   -8.001000E+3   -8.001000E+3   8.999955E+1   -8.001000E+3   -8.001000E+3   -4.020808E-1   -1.278065E-2   -2.321012E-4   3.076932E-4   -3.076950E-4   -2.320988E-4   3.854168E-4   1.270282E+2   2.170278E+2   
1.971310E+3   2.151751E+1   2.151751E+1   -8.502000E+3   -8.502000E+3   8.999955E+1   -8.501000E+3   -8.501000E+3   -3.601245E-1   -3.134987E-3   -2.133901E-4   2.700479E-4   -2.700496E-4   -2.133879E-4   3.441819E-4   1.283156E+2   2.183151E+2   
1.995601E+3   2.151919E+1   2.151919E+1   -9.001000E+3   -9.001000E+3   8.999955E+1   -9.001000E+3   -9.001000E+3   -3.206546E-1   4.402881E-3   -1.947697E-4   2.356571E-4   -2.356586E-4   -1.947679E-4   3.057279E-4   1.295736E+2   2.195732E+2   
2.019895E+3   2.151629E+1   2.151629E+1   -9.502000E+3   -9.502000E+3   8.999955E+1   -9.501000E+3   -9.501000E+3   -2.740219E-1   2.757191E-3   -1.657782E-4   2.020554E-4   -2.020567E-4   -1.657766E-4   2.613596E-4   1.293675E+2   2.193670E+2   
2.044193E+3   2.151290E+1   2.151290E+1   -1.000100E+4   -1.000100E+4   8.999955E+1   -1.000100E+4   -1.000100E+4   -2.316989E-1   -2.646492E-3   -1.368749E-4   1.741643E-4   -1.741654E-4   -1.368736E-4   2.215129E-4   1.281636E+2   2.181632E+2   
2.068134E+3   2.150121E+1   2.150121E+1   -1.050200E+4   -1.050200E+4   8.999955E+1   -1.050100E+4   -1.050100E+4   -1.910518E-1   -1.470695E-2   -1.045631E-4   1.519554E-4   -1.519563E-4   -1.045619E-4   1.844557E-4   1.245325E+2   2.145321E+2   
2.092162E+3   2.147549E+1   2.147549E+1   -1.100200E+4   -1.100200E+4   8.999955E+1   -1.100200E+4   -1.100200E+4   -1.494991E-1   -3.282564E-2   -6.769483E-5   1.331092E-4   -1.331097E-4   -6.769379E-5   1.493340E-4   1.169564E+2   2.069559E+2   
2.116644E+3   2.148101E+1   2.148101E+1   -1.150200E+4   -1.150200E+4   8.999955E+1   -1.150100E+4   -1.150100E+4   -1.130662E-1   -5.351681E-2   -3.218517E-5   1.197864E-4   -1.197867E-4   -3.218423E-5   1.240350E-4   1.050395E+2   1.950390E+2   
2.141146E+3   2.146511E+1   2.146511E+1   -1.200200E+4   -1.200200E+4   8.999955E+1   -1.200100E+4   -1.200100E+4   -7.825875E-2   -7.613422E-2   3.628477E-6   1.089565E-4   -1.089564E-4   3.629332E-6   1.090169E-4   8.809264E+1   1.780922E+2   
2.165577E+3   2.144769E+1   2.144769E+1   -1.250200E+4   -1.250200E+4   8.999955E+1   -1.250200E+4   -1.250200E+4   -4.122013E-2   -1.054485E-1   4.521486E-5   1.009283E-4   -1.009280E-4   4.521565E-5   1.105935E-4   6.586811E+1   1.558677E+2   
2.189486E+3   2.138040E+1   2.138040E+1   -1.300200E+4   -1.300200E+4   8.999955E+1   -1.300200E+4   -1.300200E+4   -1.152305E-2   -1.305599E-1   7.962354E-5   9.556254E-5   -9.556191E-5   7.962429E-5   1.243869E-4   5.019864E+1   1.401982E+2   
2.213978E+3   2.137789E+1   2.137789E+1   -1.350200E+4   -1.350200E+4   8.999955E+1   -1.350100E+4   -1.350100E+4   2.159992E-2   -1.587611E-1   1.181296E-4   8.970633E-5   -8.970540E-5   1.181303E-4   1.483301E-4   3.721265E+1   1.272122E+2   
2.238494E+3   2.136099E+1   2.136099E+1   -1.400100E+4   -1.400100E+4   8.999955E+1   -1.400100E+4   -1.400100E+4   5.711458E-2   -1.912172E-1   1.608861E-4   8.490545E-5   -8.490419E-5   1.608868E-4   1.819156E-4   2.782224E+1   1.178218E+2   
2.262476E+3   2.132549E+1   2.132549E+1   -1.450200E+4   -1.450200E+4   8.999955E+1   -1.450200E+4   -1.450200E+4   8.806012E-2   -2.205093E-1   1.988122E-4   8.139624E-5   -8.139468E-5   1.988129E-4   2.148294E-4   2.226481E+1   1.122644E+2   
2.286407E+3   2.135439E+1   2.135439E+1   -1.500200E+4   -1.500200E+4   8.999955E+1   -1.500200E+4   -1.500200E+4   1.169986E-1   -2.495491E-1   2.353713E-4   7.921234E-5   -7.921049E-5   2.353719E-4   2.483430E-4   1.860025E+1   1.085998E+2   
2.310911E+3   2.135989E+1   2.135989E+1   -1.550200E+4   -1.550200E+4   8.999955E+1   -1.550100E+4   -1.550100E+4   1.488522E-1   -2.803477E-1   2.750322E-4   7.603119E-5   -7.602903E-5   2.750328E-4   2.853479E-4   1.545318E+1   1.054527E+2   
2.335951E+3   2.136740E+1   2.136740E+1   -1.600100E+4   -1.600100E+4   8.999955E+1   -1.600100E+4   -1.600100E+4   1.819152E-1   -3.143808E-1   3.176189E-4   7.410522E-5   -7.410272E-5   3.176194E-4   3.261492E-4   1.313302E+1   1.031326E+2   
2.360905E+3   2.136440E+1   2.136440E+1   -1.650200E+4   -1.650200E+4   8.999955E+1   -1.650200E+4   -1.650200E+4   2.129251E-1   -3.481768E-1   3.587523E-4   7.354892E-5   -7.354610E-5   3.587529E-4   3.662140E-4   1.158585E+1   1.015854E+2   
2.386453E+3   2.136459E+1   2.136459E+1   -1.700200E+4   -1.700200E+4   8.999955E+1   -1.700200E+4   -1.700200E+4   2.458349E-1   -3.818595E-1   4.009763E-4   7.150349E-5   -7.150034E-5   4.009768E-4   4.073017E-4   1.011090E+1   1.001105E+2   
2.412448E+3   2.134789E+1   2.134789E+1   -1.750200E+4   -1.750200E+4   8.999955E+1   -1.750200E+4   -1.750200E+4   2.714578E-1   -4.109825E-1   4.357574E-4   7.184200E-5   -7.183858E-5   4.357580E-4   4.416399E-4   9.361964E+0   9.936151E+1   
2.438955E+3   2.134490E+1   2.134490E+1   -1.800200E+4   -1.800200E+4   8.999955E+1   -1.800200E+4   -1.800200E+4   3.039138E-1   -4.443879E-1   4.774091E-4   6.994946E-5   -6.994571E-5   4.774097E-4   4.825064E-4   8.335603E+0   9.833515E+1   
2.465451E+3   2.134661E+1   2.134661E+1   -1.850200E+4   -1.850200E+4   8.999955E+1   -1.850200E+4   -1.850200E+4   3.352628E-1   -4.777237E-1   5.184383E-4   6.883434E-5   -6.883027E-5   5.184388E-4   5.229880E-4   7.563068E+0   9.756262E+1   
2.492484E+3   2.136270E+1   2.136270E+1   -1.900300E+4   -1.900300E+4   8.999955E+1   -1.900200E+4   -1.900200E+4   3.622568E-1   -5.096107E-1   5.558115E-4   6.999427E-5   -6.998991E-5   5.558120E-4   5.602014E-4   7.177571E+0   9.717712E+1   
2.519447E+3   2.133679E+1   2.133679E+1   -1.950200E+4   -1.950200E+4   8.999955E+1   -1.950200E+4   -1.950200E+4   3.905710E-1   -5.411928E-1   5.938805E-4   6.996867E-5   -6.996400E-5   5.938811E-4   5.979881E-4   6.719388E+0   9.671894E+1   
2.547484E+3   2.131521E+1   2.131521E+1   -2.000100E+4   -2.000100E+4   8.999955E+1   -2.000100E+4   -2.000100E+4   4.188395E-1   -5.725277E-1   6.315448E-4   6.981250E-5   -6.980754E-5   6.315453E-4   6.353917E-4   6.308005E+0   9.630755E+1   
2.590176E+3   2.134319E+1   2.134319E+1   -1.950200E+4   -1.950200E+4   8.999955E+1   -1.950200E+4   -1.950200E+4   3.919916E-1   -5.438373E-1   5.964898E-4   7.067367E-5   -7.066899E-5   5.964904E-4   6.006620E-4   6.757052E+0   9.675660E+1   
2.619931E+3   2.133889E+1   2.133889E+1   -1.900200E+4   -1.900200E+4   8.999955E+1   -1.900200E+4   -1.900200E+4   3.637667E-1   -5.107119E-1   5.574486E-4   6.960450E-5   -6.960012E-5   5.574492E-4   5.617773E-4   7.117267E+0   9.711682E+1   
2.649178E+3   2.134271E+1   2.134271E+1   -1.850200E+4   -1.850200E+4   8.999955E+1   -1.850200E+4   -1.850200E+4   3.300471E-1   -4.762570E-1   5.143356E-4   7.173800E-5   -7.173396E-5   5.143362E-4   5.193144E-4   7.940220E+0   9.793977E+1   
2.677678E+3   2.133981E+1   2.133981E+1   -1.800200E+4   -1.800200E+4   8.999955E+1   -1.800200E+4   -1.800200E+4   2.971175E-1   -4.413017E-1   4.712837E-4   7.295022E-5   -7.294652E-5   4.712843E-4   4.768963E-4   8.799008E+0   9.879856E+1   
2.705642E+3   2.134039E+1   2.134039E+1   -1.750200E+4   -1.750200E+4   8.999955E+1   -1.750200E+4   -1.750200E+4   2.723834E-1   -4.127608E-1   4.374937E-4   7.233817E-5   -7.233473E-5   4.374942E-4   4.434338E-4   9.388726E+0   9.938828E+1   
2.733588E+3   2.136590E+1   2.136590E+1   -1.700200E+4   -1.700200E+4   8.999955E+1   -1.700200E+4   -1.700200E+4   2.411855E-1   -3.805356E-1   3.973095E-4   7.408086E-5   -7.407774E-5   3.973100E-4   4.041569E-4   1.056188E+1   1.005614E+2   
2.761938E+3   2.136682E+1   2.136682E+1   -1.650200E+4   -1.650200E+4   8.999955E+1   -1.650200E+4   -1.650200E+4   2.153952E-1   -3.505174E-1   3.617866E-4   7.327046E-5   -7.326762E-5   3.617872E-4   3.691316E-4   1.144891E+1   1.014485E+2   
2.789393E+3   2.138519E+1   2.138519E+1   -1.600100E+4   -1.600100E+4   8.999955E+1   -1.600100E+4   -1.600100E+4   1.803905E-1   -3.154846E-1   3.174378E-4   7.597510E-5   -7.597261E-5   3.174384E-4   3.264031E-4   1.345989E+1   1.034594E+2   
2.816797E+3   2.139568E+1   2.139568E+1   -1.550200E+4   -1.550200E+4   8.999955E+1   -1.550100E+4   -1.550100E+4   1.499122E-1   -2.853108E-1   2.789580E-4   7.854919E-5   -7.854700E-5   2.789586E-4   2.898060E-4   1.572620E+1   1.057257E+2   
2.843748E+3   2.142660E+1   2.142660E+1   -1.500200E+4   -1.500200E+4   8.999955E+1   -1.500100E+4   -1.500100E+4   1.201863E-1   -2.536469E-1   2.399936E-4   7.957069E-5   -7.956880E-5   2.399942E-4   2.528407E-4   1.834312E+1   1.083427E+2   
2.870771E+3   2.141360E+1   2.141360E+1   -1.450200E+4   -1.450200E+4   8.999955E+1   -1.450200E+4   -1.450200E+4   8.573480E-2   -2.210750E-1   1.977958E-4   8.350336E-5   -8.350181E-5   1.977965E-4   2.146998E-4   2.288799E+1   1.128875E+2   
2.896632E+3   2.140289E+1   2.140289E+1   -1.400100E+4   -1.400100E+4   8.999955E+1   -1.400100E+4   -1.400100E+4   5.393578E-2   -1.897659E-1   1.580225E-4   8.630378E-5   -8.630254E-5   1.580232E-4   1.800540E-4   2.864110E+1   1.186407E+2   
2.922041E+3   2.146929E+1   2.146929E+1   -1.350200E+4   -1.350200E+4   8.999955E+1   -1.350100E+4   -1.350100E+4   2.156711E-2   -1.598404E-1   1.188251E-4   9.044986E-5   -9.044893E-5   1.188258E-4   1.493338E-4   3.727844E+1   1.272780E+2   
2.948839E+3   2.147979E+1   2.147979E+1   -1.300200E+4   -1.300200E+4   8.999955E+1   -1.300200E+4   -1.300200E+4   -9.885732E-3   -1.321283E-1   8.164254E-5   9.538928E-5   -9.538864E-5   8.164329E-5   1.255572E-4   4.944018E+1   1.394397E+2   
2.974331E+3   2.155959E+1   2.155959E+1   -1.250200E+4   -1.250200E+4   8.999955E+1   -1.250100E+4   -1.250100E+4   -4.811440E-2   -1.033684E-1   3.971149E-5   1.046723E-4   -1.046719E-4   3.971232E-5   1.119522E-4   6.922381E+1   1.592234E+2   
2.999755E+3   2.161089E+1   2.161089E+1   -1.200100E+4   -1.200100E+4   8.999955E+1   -1.200100E+4   -1.200100E+4   -7.784813E-2   -7.717170E-2   4.561657E-6   1.093422E-4   -1.093421E-4   4.562516E-6   1.094373E-4   8.761106E+1   1.776106E+2   
3.025302E+3   2.164239E+1   2.164239E+1   -1.150200E+4   -1.150200E+4   8.999955E+1   -1.150100E+4   -1.150100E+4   -1.146186E-1   -5.219102E-2   -3.399252E-5   1.200581E-4   -1.200584E-4   -3.399157E-5   1.247776E-4   1.058086E+2   1.958082E+2   
3.052051E+3   2.167211E+1   2.167211E+1   -1.100200E+4   -1.100200E+4   8.999955E+1   -1.100200E+4   -1.100200E+4   -1.511924E-1   -3.428788E-2   -6.773898E-5   1.353434E-4   -1.353439E-4   -6.773792E-5   1.513486E-4   1.165878E+2   2.065874E+2   
3.078048E+3   2.167281E+1   2.167281E+1   -1.050200E+4   -1.050200E+4   8.999955E+1   -1.050100E+4   -1.050100E+4   -1.867538E-1   -1.784194E-2   -9.991410E-5   1.508462E-4   -1.508470E-4   -9.991292E-5   1.809348E-4   1.235188E+2   2.135183E+2   
3.103959E+3   2.169799E+1   2.169799E+1   -1.000100E+4   -1.000100E+4   8.999955E+1   -1.000000E+4   -1.000000E+4   -2.314376E-1   -3.201278E-3   -1.363510E-4   1.743396E-4   -1.743406E-4   -1.363496E-4   2.213275E-4   1.280290E+2   2.180285E+2   
3.129146E+3   2.174069E+1   2.174069E+1   -9.501000E+3   -9.501000E+3   8.999955E+1   -9.501000E+3   -9.501000E+3   -2.721568E-1   1.674654E-3   -1.639449E-4   2.013889E-4   -2.013902E-4   -1.639433E-4   2.596833E-4   1.291480E+2   2.191476E+2   
3.154299E+3   2.176501E+1   2.176501E+1   -9.001000E+3   -9.001000E+3   8.999955E+1   -9.001000E+3   -9.001000E+3   -3.175917E-1   1.610295E-3   -1.910866E-4   2.352387E-4   -2.352402E-4   -1.910848E-4   3.030699E-4   1.290873E+2   2.190868E+2   
3.179995E+3   2.178671E+1   2.178671E+1   -8.502000E+3   -8.502000E+3   8.999955E+1   -8.501000E+3   -8.501000E+3   -3.569825E-1   -5.764102E-3   -2.097679E-4   2.694617E-4   -2.694634E-4   -2.097658E-4   3.414853E-4   1.278997E+2   2.178992E+2   
3.205188E+3   2.180419E+1   2.180419E+1   -8.001000E+3   -8.001000E+3   8.999955E+1   -8.000000E+3   -8.000000E+3   -3.984983E-1   -1.567815E-2   -2.280376E-4   3.069580E-4   -3.069598E-4   -2.280352E-4   3.823930E-4   1.266085E+2   2.166080E+2   
3.231332E+3   2.184490E+1   2.184490E+1   -7.501000E+3   -7.501000E+3   8.999955E+1   -7.501000E+3   -7.501000E+3   -4.375936E-1   -2.767683E-2   -2.434778E-4   3.440422E-4   -3.440441E-4   -2.434751E-4   4.214813E-4   1.252869E+2   2.152865E+2   
3.257849E+3   2.186840E+1   2.186840E+1   -7.002000E+3   -7.002000E+3   8.999955E+1   -7.001000E+3   -7.001000E+3   -4.728863E-1   -3.962654E-2   -2.566752E-4   3.782644E-4   -3.782664E-4   -2.566722E-4   4.571281E-4   1.241593E+2   2.141588E+2   
3.283935E+3   2.188979E+1   2.188979E+1   -6.502000E+3   -6.502000E+3   8.999955E+1   -6.501000E+3   -6.501000E+3   -5.025053E-1   -5.611252E-2   -2.634719E-4   4.112873E-4   -4.112893E-4   -2.634687E-4   4.884410E-4   1.226438E+2   2.126433E+2   
3.309082E+3   2.192620E+1   2.192620E+1   -6.001000E+3   -6.001000E+3   8.999955E+1   -6.001000E+3   -6.001000E+3   -5.342336E-1   -6.876180E-2   -2.740731E-4   4.433233E-4   -4.433255E-4   -2.740696E-4   5.212021E-4   1.217254E+2   2.117249E+2   
3.335240E+3   2.194381E+1   2.194381E+1   -5.501000E+3   -5.501000E+3   8.999955E+1   -5.501000E+3   -5.501000E+3   -5.595862E-1   -8.105838E-2   -2.810934E-4   4.703804E-4   -4.703826E-4   -2.810897E-4   5.479701E-4   1.208620E+2   2.108616E+2   
3.361691E+3   2.197030E+1   2.197030E+1   -5.002000E+3   -5.002000E+3   8.999955E+1   -5.001000E+3   -5.001000E+3   -5.848295E-1   -9.473169E-2   -2.871359E-4   4.982734E-4   -4.982757E-4   -2.871320E-4   5.750856E-4   1.199532E+2   2.099528E+2   
3.397237E+3   2.198062E+1   2.198062E+1   -4.801000E+3   -4.801000E+3   8.999955E+1   -4.801000E+3   -4.801000E+3   -5.937690E-1   -9.980023E-2   -2.891258E-4   5.083021E-4   -5.083044E-4   -2.891218E-4   5.847776E-4   1.196315E+2   2.096311E+2   
3.421989E+3   2.202450E+1   2.202450E+1   -4.601000E+3   -4.601000E+3   8.999955E+1   -4.601000E+3   -4.601000E+3   -6.037948E-1   -1.041775E-1   -2.922237E-4   5.186785E-4   -5.186808E-4   -2.922196E-4   5.953335E-4   1.193969E+2   2.093965E+2   
3.446221E+3   2.203961E+1   2.203961E+1   -4.401000E+3   -4.401000E+3   8.999955E+1   -4.401000E+3   -4.401000E+3   -6.128770E-1   -1.093166E-1   -2.942521E-4   5.288603E-4   -5.288627E-4   -2.942480E-4   6.052087E-4   1.190911E+2   2.090906E+2   
3.469935E+3   2.204690E+1   2.204690E+1   -4.201000E+3   -4.201000E+3   8.999955E+1   -4.201000E+3   -4.201000E+3   -6.190424E-1   -1.140870E-1   -2.947798E-4   5.366263E-4   -5.366286E-4   -2.947756E-4   6.122605E-4   1.187809E+2   2.087804E+2   
3.494114E+3   2.206759E+1   2.206759E+1   -4.000000E+3   -4.000000E+3   8.999955E+1   -4.000000E+3   -4.000000E+3   -6.253801E-1   -1.200583E-1   -2.946148E-4   5.453205E-4   -5.453228E-4   -2.946105E-4   6.198163E-4   1.183806E+2   2.083801E+2   
3.517764E+3   2.207839E+1   2.207839E+1   -3.800000E+3   -3.800000E+3   8.999955E+1   -3.800000E+3   -3.800000E+3   -6.333614E-1   -1.248067E-1   -2.962434E-4   5.544229E-4   -5.544253E-4   -2.962390E-4   6.286056E-4   1.181168E+2   2.081164E+2   
3.541043E+3   2.209670E+1   2.209670E+1   -3.601000E+3   -3.601000E+3   8.999955E+1   -3.600000E+3   -3.600000E+3   -6.394786E-1   -1.302040E-1   -2.963269E-4   5.625706E-4   -5.625730E-4   -2.963225E-4   6.358422E-4   1.177774E+2   2.077770E+2   
3.565243E+3   2.210790E+1   2.210790E+1   -3.401000E+3   -3.401000E+3   8.999955E+1   -3.401000E+3   -3.401000E+3   -6.472713E-1   -1.353862E-1   -2.975552E-4   5.718218E-4   -5.718241E-4   -2.975507E-4   6.446078E-4   1.174908E+2   2.074904E+2   
3.589030E+3   2.211239E+1   2.211239E+1   -3.201000E+3   -3.201000E+3   8.999955E+1   -3.201000E+3   -3.201000E+3   -6.537621E-1   -1.385630E-1   -2.993336E-4   5.787680E-4   -5.787703E-4   -2.993290E-4   6.515926E-4   1.173476E+2   2.073471E+2   
3.612728E+3   2.213430E+1   2.213430E+1   -3.001000E+3   -3.001000E+3   8.999955E+1   -3.001000E+3   -3.001000E+3   -6.608453E-1   -1.443754E-1   -2.997199E-4   5.879111E-4   -5.879134E-4   -2.997153E-4   6.599026E-4   1.170127E+2   2.070123E+2   
3.636926E+3   2.214269E+1   2.214269E+1   -2.801000E+3   -2.801000E+3   8.999955E+1   -2.801000E+3   -2.801000E+3   -6.668239E-1   -1.489005E-1   -3.002983E-4   5.953745E-4   -5.953769E-4   -3.002936E-4   6.668207E-4   1.167657E+2   2.067653E+2   
3.661141E+3   2.215750E+1   2.215750E+1   -2.601000E+3   -2.601000E+3   8.999955E+1   -2.601000E+3   -2.601000E+3   -6.746533E-1   -1.538543E-1   -3.017001E-4   6.045008E-4   -6.045032E-4   -3.016953E-4   6.756065E-4   1.165233E+2   2.065229E+2   
3.684880E+3   2.217001E+1   2.217001E+1   -2.401000E+3   -2.401000E+3   8.999955E+1   -2.401000E+3   -2.401000E+3   -6.815745E-1   -1.591060E-1   -3.023609E-4   6.131498E-4   -6.131522E-4   -3.023561E-4   6.836482E-4   1.162492E+2   2.062487E+2   
3.709073E+3   2.218090E+1   2.218090E+1   -2.201000E+3   -2.201000E+3   8.999955E+1   -2.200000E+3   -2.200000E+3   -6.869255E-1   -1.640199E-1   -3.023062E-4   6.204053E-4   -6.204076E-4   -3.023013E-4   6.901389E-4   1.159787E+2   2.059782E+2   
3.732806E+3   2.218591E+1   2.218591E+1   -2.000000E+3   -2.000000E+3   8.999955E+1   -2.000000E+3   -2.000000E+3   -6.899258E-1   -1.693772E-1   -3.005512E-4   6.262072E-4   -6.262095E-4   -3.005463E-4   6.945981E-4   1.156389E+2   2.056385E+2   
3.756094E+3   2.218191E+1   2.218191E+1   -1.800000E+3   -1.800000E+3   8.999955E+1   -1.800000E+3   -1.800000E+3   -6.976151E-1   -1.760024E-1   -3.007615E-4   6.363427E-4   -6.363451E-4   -3.007565E-4   7.038391E-4   1.152973E+2   2.052969E+2   
3.779834E+3   2.220001E+1   2.220001E+1   -1.601000E+3   -1.601000E+3   8.999955E+1   -1.601000E+3   -1.601000E+3   -7.041771E-1   -1.792732E-1   -3.025202E-4   6.434046E-4   -6.434070E-4   -3.025152E-4   7.109768E-4   1.151823E+2   2.051818E+2   
3.804080E+3   2.220321E+1   2.220321E+1   -1.401000E+3   -1.401000E+3   8.999955E+1   -1.401000E+3   -1.401000E+3   -7.094662E-1   -1.853359E-1   -3.016672E-4   6.513795E-4   -6.513818E-4   -3.016621E-4   7.178428E-4   1.148498E+2   2.048494E+2   
3.827834E+3   2.220931E+1   2.220931E+1   -1.201000E+3   -1.201000E+3   8.999955E+1   -1.201000E+3   -1.201000E+3   -7.165652E-1   -1.927502E-1   -3.010014E-4   6.616016E-4   -6.616040E-4   -3.009962E-4   7.268552E-4   1.144636E+2   2.044631E+2   
3.852845E+3   2.222680E+1   2.222680E+1   -1.002000E+3   -1.002000E+3   8.999955E+1   -1.001000E+3   -1.001000E+3   -7.232386E-1   -1.995368E-1   -3.004969E-4   6.710889E-4   -6.710912E-4   -3.004916E-4   7.352950E-4   1.141216E+2   2.041212E+2   
3.876884E+3   2.223419E+1   2.223419E+1   -8.020000E+2   -8.020000E+2   8.999955E+1   -8.010000E+2   -8.010000E+2   -7.292369E-1   -2.088351E-1   -2.979241E-4   6.817472E-4   -6.817495E-4   -2.979187E-4   7.440014E-4   1.136054E+2   2.036049E+2   
3.900873E+3   2.224249E+1   2.224249E+1   -6.010000E+2   -6.010000E+2   8.999955E+1   -6.010000E+2   -6.010000E+2   -7.400545E-1   -2.209708E-1   -2.963545E-4   6.978820E-4   -6.978843E-4   -2.963490E-4   7.581987E-4   1.130084E+2   2.030080E+2   
3.924406E+3   2.223580E+1   2.223580E+1   -4.010000E+2   -4.010000E+2   8.999955E+1   -4.010000E+2   -4.010000E+2   -7.503721E-1   -2.344844E-1   -2.935726E-4   7.145628E-4   -7.145651E-4   -2.935669E-4   7.725185E-4   1.123349E+2   2.023345E+2   
3.947988E+3   2.222961E+1   2.222961E+1   -2.010000E+2   -2.010000E+2   8.999955E+1   -2.010000E+2   -2.010000E+2   -7.643367E-1   -2.513860E-1   -2.907276E-4   7.362145E-4   -7.362168E-4   -2.907218E-4   7.915393E-4   1.115488E+2   2.015484E+2   
3.971065E+3   2.224261E+1   2.224261E+1   -1.000000E+0   -1.000000E+0   8.999955E+1   0.000000E+0   0.000000E+0   -7.502472E-1   -2.503253E-1   -2.830006E-4   7.250242E-4   -7.250264E-4   -2.829949E-4   7.782991E-4   1.113223E+2   2.013219E+2   
4.007902E+3   2.224951E+1   2.224951E+1   1.970000E+2   1.970000E+2   8.999955E+1   1.970000E+2   1.970000E+2   -3.777681E-1   3.337978E-2   -2.481437E-4   2.588473E-4   -2.588492E-4   -2.481416E-4   3.585766E-4   1.337906E+2   2.237901E+2   
4.033142E+3   2.224740E+1   2.224740E+1   3.970000E+2   3.970000E+2   8.999955E+1   3.970000E+2   3.970000E+2   1.744887E-1   2.415576E-1   -5.567365E-5   -2.907758E-4   2.907753E-4   -5.567593E-5   2.960576E-4   -1.008390E+2   -1.083946E+1   
4.058827E+3   2.224761E+1   2.224761E+1   5.960000E+2   5.960000E+2   8.999955E+1   5.970000E+2   5.970000E+2   3.914274E-1   1.809819E-1   1.142654E-4   -4.118342E-4   4.118351E-4   1.142621E-4   4.273921E-4   -7.449307E+1   1.550648E+1   
4.084070E+3   2.222610E+1   2.222610E+1   7.960000E+2   7.960000E+2   8.999955E+1   7.960000E+2   7.960000E+2   5.376558E-1   1.862054E-1   1.982944E-4   -5.241192E-4   5.241207E-4   1.982903E-4   5.603763E-4   -6.927644E+1   2.072311E+1   
4.109757E+3   2.224551E+1   2.224551E+1   9.960000E+2   9.960000E+2   8.999955E+1   9.970000E+2   9.970000E+2   6.416089E-1   1.880693E-1   2.592559E-4   -6.027098E-4   6.027118E-4   2.592512E-4   6.561042E-4   -6.672502E+1   2.327453E+1   
4.135294E+3   2.223531E+1   2.223531E+1   1.197000E+3   1.197000E+3   8.999955E+1   1.197000E+3   1.197000E+3   6.987489E-1   1.666516E-1   3.076364E-4   -6.309562E-4   6.309586E-4   3.076314E-4   7.019586E-4   -6.400745E+1   2.599210E+1   
4.160791E+3   2.223010E+1   2.223010E+1   1.397000E+3   1.397000E+3   8.999955E+1   1.397000E+3   1.397000E+3   7.086983E-1   1.592940E-1   3.184649E-4   -6.334571E-4   6.334596E-4   3.184600E-4   7.090048E-4   -6.330944E+1   2.669011E+1   
4.186187E+3   2.223708E+1   2.223708E+1   1.597000E+3   1.597000E+3   8.999955E+1   1.597000E+3   1.597000E+3   7.085477E-1   1.570182E-1   3.198829E-4   -6.318287E-4   6.318312E-4   3.198779E-4   7.081896E-4   -6.314777E+1   2.685178E+1   
4.212244E+3   2.222430E+1   2.222430E+1   1.797000E+3   1.797000E+3   8.999955E+1   1.798000E+3   1.798000E+3   7.061137E-1   1.534462E-1   3.207936E-4   -6.276377E-4   6.276402E-4   3.207887E-4   7.048671E-4   -6.292785E+1   2.707170E+1   
4.237691E+3   2.222949E+1   2.222949E+1   1.997000E+3   1.997000E+3   8.999955E+1   1.998000E+3   1.998000E+3   7.022726E-1   1.484120E-1   3.218315E-4   -6.214255E-4   6.214280E-4   3.218266E-4   6.998180E-4   -6.262071E+1   2.737884E+1   
4.275945E+3   2.220391E+1   2.220391E+1   2.497000E+3   2.497000E+3   8.999955E+1   2.497000E+3   2.497000E+3   6.895260E-1   1.379200E-1   3.211577E-4   -6.049506E-4   6.049531E-4   3.211529E-4   6.849142E-4   -6.203695E+1   2.796260E+1   
4.302889E+3   2.221160E+1   2.221160E+1   2.997000E+3   2.997000E+3   8.999955E+1   2.997000E+3   2.997000E+3   6.759493E-1   1.263443E-1   3.207054E-4   -5.871359E-4   5.871384E-4   3.207008E-4   6.690146E-4   -6.135575E+1   2.864380E+1   
4.329824E+3   2.220989E+1   2.220989E+1   3.497000E+3   3.497000E+3   8.999955E+1   3.497000E+3   3.497000E+3   6.590176E-1   1.174478E-1   3.164704E-4   -5.686100E-4   5.686125E-4   3.164659E-4   6.507463E-4   -6.090107E+1   2.909848E+1   
4.356434E+3   2.221481E+1   2.221481E+1   3.997000E+3   3.997000E+3   8.999955E+1   3.998000E+3   3.998000E+3   6.418272E-1   1.044728E-1   3.147833E-4   -5.471742E-4   5.471767E-4   3.147790E-4   6.312592E-4   -6.008866E+1   2.991089E+1   
4.383418E+3   2.219631E+1   2.219631E+1   4.497000E+3   4.497000E+3   8.999955E+1   4.497000E+3   4.497000E+3   6.210106E-1   9.157286E-2   3.108768E-4   -5.230902E-4   5.230926E-4   3.108727E-4   6.084963E-4   -5.927663E+1   3.072292E+1   
4.410410E+3   2.219311E+1   2.219311E+1   4.996000E+3   4.996000E+3   8.999955E+1   4.997000E+3   4.997000E+3   5.979066E-1   7.802898E-2   3.060285E-4   -4.968752E-4   4.968776E-4   3.060246E-4   5.835567E-4   -5.837083E+1   3.162872E+1   
4.437317E+3   2.218371E+1   2.218371E+1   5.497000E+3   5.497000E+3   8.999955E+1   5.497000E+3   5.497000E+3   5.726428E-1   6.602330E-2   2.988686E-4   -4.700780E-4   4.700804E-4   2.988649E-4   5.570420E-4   -5.755241E+1   3.244714E+1   
4.464261E+3   2.218499E+1   2.218499E+1   5.997000E+3   5.997000E+3   8.999955E+1   5.997000E+3   5.997000E+3   5.449044E-1   5.380134E-2   2.903714E-4   -4.412954E-4   4.412977E-4   2.903679E-4   5.282586E-4   -5.665517E+1   3.334438E+1   
4.491183E+3   2.215649E+1   2.215649E+1   6.496000E+3   6.496000E+3   8.999955E+1   6.497000E+3   6.497000E+3   5.191797E-1   3.774531E-2   2.856198E-4   -4.114567E-4   4.114589E-4   2.856166E-4   5.008745E-4   -5.523288E+1   3.476667E+1   
4.517626E+3   2.215331E+1   2.215331E+1   6.996000E+3   6.996000E+3   8.999955E+1   6.996000E+3   6.996000E+3   4.853685E-1   2.364788E-2   2.747320E-4   -3.769059E-4   3.769080E-4   2.747290E-4   4.664072E-4   -5.391116E+1   3.608839E+1   
4.544440E+3   2.213751E+1   2.213751E+1   7.497000E+3   7.497000E+3   8.999955E+1   7.497000E+3   7.497000E+3   4.496191E-1   1.084663E-2   2.618257E-4   -3.417766E-4   3.417786E-4   2.618230E-4   4.305391E-4   -5.254526E+1   3.745429E+1   
4.570875E+3   2.213690E+1   2.213690E+1   7.997000E+3   7.997000E+3   8.999955E+1   7.998000E+3   7.998000E+3   4.110502E-1   -1.659206E-3   2.470366E-4   -3.047461E-4   3.047481E-4   2.470342E-4   3.922974E-4   -5.097072E+1   3.902883E+1   
4.597863E+3   2.212771E+1   2.212771E+1   8.496000E+3   8.496000E+3   8.999955E+1   8.497000E+3   8.497000E+3   3.717711E-1   -1.291838E-2   2.309964E-4   -2.680179E-4   2.680197E-4   2.309943E-4   3.538261E-4   -4.924296E+1   4.075659E+1   
4.624774E+3   2.211111E+1   2.211111E+1   8.996000E+3   8.996000E+3   8.999955E+1   8.997000E+3   8.997000E+3   3.276229E-1   -1.706189E-2   2.073277E-4   -2.324077E-4   2.324093E-4   2.073259E-4   3.114452E-4   -4.826428E+1   4.173527E+1   
4.652177E+3   2.209438E+1   2.209438E+1   9.497000E+3   9.497000E+3   8.999955E+1   9.497000E+3   9.497000E+3   2.849098E-1   -1.869535E-2   1.828543E-4   -1.995377E-4   1.995391E-4   1.828527E-4   2.706492E-4   -4.749817E+1   4.250138E+1   
4.678582E+3   2.208041E+1   2.208041E+1   9.997000E+3   9.997000E+3   8.999955E+1   9.998000E+3   9.998000E+3   2.427675E-1   -1.126947E-2   1.527191E-4   -1.731284E-4   1.731296E-4   1.527178E-4   2.308605E-4   -4.858400E+1   4.141555E+1   
4.705861E+3   2.207079E+1   2.207079E+1   1.049700E+4   1.049700E+4   8.999955E+1   1.049700E+4   1.049700E+4   2.029485E-1   -9.454525E-4   1.220534E-4   -1.503787E-4   1.503797E-4   1.220523E-4   1.936771E-4   -5.093582E+1   3.906373E+1   
4.733099E+3   2.206170E+1   2.206170E+1   1.099600E+4   1.099600E+4   8.999955E+1   1.099700E+4   1.099700E+4   1.628254E-1   1.618209E-2   8.669733E-5   -1.319358E-4   1.319365E-4   8.669630E-5   1.578717E-4   -5.669038E+1   3.330917E+1   
4.759954E+3   2.205111E+1   2.205111E+1   1.149700E+4   1.149700E+4   8.999955E+1   1.149700E+4   1.149700E+4   1.265277E-1   3.926228E-2   4.968542E-5   -1.203054E-4   1.203058E-4   4.968447E-5   1.301615E-4   -6.755966E+1   2.243989E+1   
4.787248E+3   2.202300E+1   2.202300E+1   1.199700E+4   1.199700E+4   8.999955E+1   1.199700E+4   1.199700E+4   8.763282E-2   6.425790E-2   9.850235E-6   -1.080186E-4   1.080187E-4   9.849386E-6   1.084668E-4   -8.478960E+1   5.209951E+0   
4.814073E+3   2.201699E+1   2.201699E+1   1.249600E+4   1.249600E+4   8.999955E+1   1.249700E+4   1.249700E+4   5.900676E-2   8.765592E-2   -2.278228E-5   -1.023082E-4   1.023080E-4   -2.278308E-5   1.048141E-4   -1.025540E+2   -1.255441E+1   
4.841415E+3   2.193539E+1   2.193539E+1   1.299600E+4   1.299600E+4   8.999955E+1   1.299600E+4   1.299600E+4   2.497692E-2   1.166491E-1   -6.235570E-5   -9.630487E-5   9.630438E-5   -6.235646E-5   1.147295E-4   -1.229223E+2   -3.292279E+1   
4.868764E+3   2.194521E+1   2.194521E+1   1.349700E+4   1.349700E+4   8.999955E+1   1.349700E+4   1.349700E+4   -1.038581E-2   1.453272E-1   -1.025178E-4   -8.909984E-5   8.909903E-5   -1.025185E-4   1.358259E-4   -1.390056E+2   -4.900603E+1   
4.895270E+3   2.190579E+1   2.190579E+1   1.399700E+4   1.399700E+4   8.999955E+1   1.399700E+4   1.399700E+4   -4.354354E-2   1.763899E-1   -1.429408E-4   -8.512426E-5   8.512313E-5   -1.429414E-4   1.663677E-4   -1.492253E+2   -5.922576E+1   
4.922616E+3   2.189559E+1   2.189559E+1   1.449600E+4   1.449600E+4   8.999955E+1   1.449700E+4   1.449700E+4   -7.005865E-2   2.033200E-1   -1.766509E-4   -8.333787E-5   8.333648E-5   -1.766515E-4   1.953221E-4   -1.547437E+2   -6.474411E+1   
4.949924E+3   2.191281E+1   2.191281E+1   1.499600E+4   1.499600E+4   8.999955E+1   1.499700E+4   1.499700E+4   -1.037120E-1   2.358057E-1   -2.183134E-4   -7.994165E-5   7.993993E-5   -2.183141E-4   2.324896E-4   -1.598884E+2   -6.988881E+1   
4.977256E+3   2.190951E+1   2.190951E+1   1.549700E+4   1.549700E+4   8.999955E+1   1.549700E+4   1.549700E+4   -1.312247E-1   2.644588E-1   -2.539399E-4   -7.856096E-5   7.855896E-5   -2.539405E-4   2.658144E-4   -1.628096E+2   -7.281004E+1   
5.004544E+3   2.190429E+1   2.190429E+1   1.599700E+4   1.599700E+4   8.999955E+1   1.599800E+4   1.599800E+4   -1.667887E-1   2.985469E-1   -2.980478E-4   -7.481073E-5   7.480839E-5   -2.980483E-4   3.072932E-4   -1.659097E+2   -7.591016E+1   
5.032829E+3   2.188760E+1   2.188760E+1   1.649600E+4   1.649600E+4   8.999955E+1   1.649700E+4   1.649700E+4   -1.924678E-1   3.297105E-1   -3.342311E-4   -7.646706E-5   7.646443E-5   -3.342317E-4   3.428668E-4   -1.671134E+2   -7.711382E+1   
5.061074E+3   2.188131E+1   2.188131E+1   1.699600E+4   1.699600E+4   8.999955E+1   1.699600E+4   1.699600E+4   -2.323039E-1   3.684874E-1   -3.839834E-4   -7.266208E-5   7.265907E-5   -3.839840E-4   3.907980E-4   -1.692845E+2   -7.928494E+1   
5.090334E+3   2.186700E+1   2.186700E+1   1.749600E+4   1.749600E+4   8.999955E+1   1.749700E+4   1.749700E+4   -2.557760E-1   3.950194E-1   -4.157497E-4   -7.287465E-5   7.287138E-5   -4.157502E-4   4.220883E-4   -1.700579E+2   -8.005837E+1   
5.119718E+3   2.186700E+1   2.186700E+1   1.799600E+4   1.799600E+4   8.999955E+1   1.799700E+4   1.799700E+4   -2.862374E-1   4.277404E-1   -4.557509E-4   -7.201026E-5   7.200668E-5   -4.557515E-4   4.614048E-4   -1.710213E+2   -8.102174E+1   
5.149013E+3   2.186569E+1   2.186569E+1   1.849600E+4   1.849600E+4   8.999955E+1   1.849600E+4   1.849600E+4   -3.166024E-1   4.619478E-1   -4.967661E-4   -7.220795E-5   7.220405E-5   -4.967667E-4   5.019866E-4   -1.717296E+2   -8.173008E+1   
5.178825E+3   2.185281E+1   2.185281E+1   1.899600E+4   1.899600E+4   8.999955E+1   1.899600E+4   1.899600E+4   -3.468598E-1   4.942745E-1   -5.363887E-4   -7.123264E-5   7.122842E-5   -5.363893E-4   5.410979E-4   -1.724354E+2   -8.243581E+1   
5.208582E+3   2.184789E+1   2.184789E+1   1.949600E+4   1.949600E+4   8.999955E+1   1.949700E+4   1.949700E+4   -3.782946E-1   5.300263E-1   -5.790959E-4   -7.166333E-5   7.165878E-5   -5.790965E-4   5.835132E-4   -1.729455E+2   -8.294594E+1   
5.239442E+3   2.183099E+1   2.183099E+1   1.999700E+4   1.999700E+4   8.999955E+1   1.999700E+4   1.999700E+4   -4.074425E-1   5.599899E-1   -6.163810E-4   -6.993904E-5   6.993420E-5   -6.163815E-4   6.203362E-4   -1.735265E+2   -8.352694E+1   
@@END Data.
@Time at end of measurement: 13:08:27
@NO Instrument  Changes.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -19502.000     -20001.000     249.500        Coercive Field: Field at which M//H changes sign
Ms  emu                                 6.315E-4       -6.661E-4      6.488E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -2.830E-4      2.851E-4       2.840E-4       Remanent Magnetization: M at H=0        
S                                       0.448          0.428          0.438          Squareness: Mr/Ms                       
S*                                      1.187          1.187          1.187          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
