@Filename: c:\vsm-lv\Will\data\AJA335e-FePtFeRh_1030nm_Tann_6\AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_90deg.VHD
@Measurement Controlfilename: C:\vsm-lv\Will\Recipes\10kOe OoP loop 90deg.VHC
@Signal Manipulation filename: c:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA335e-FePtFeRh_1030nm_Tann_6
@Date: 07 November 2019    (2019-07-11)
@Time: 12:59:55
@Test ID: AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_90deg
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 90.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Sample Temperature to 90.0977 [degC] and wait 60.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Applied Field to 9999.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 3:      Set Auto Range Signal to 13.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 5
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 5.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 10000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To: 50.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: 50.0000 [Oe] To: -50.0000 [Oe] Min Stepsize/Sweeprate =  2.0000 [Oe] Max Stepsize/Sweeprate =  2.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -50.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -10000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 4 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 50 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.706
@Y Coils Correction Factor: 0.964
@Sample Shape Correction Factor: 0.919
@Coil Angle Alpha: 42.300
@Coil Angle Beta: -47.320
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
15000.000000   1.000000
15249.000000   1.000524
15499.000000   1.000702
15750.000000   1.001233
16000.000000   1.001406
16250.000000   1.001585
16499.000000   1.001758
16749.000000   1.001937
16999.000000   1.002110
17249.000000   1.001937
17499.000000   1.002289
17749.000000   1.002289
17999.000000   1.002289
18249.000000   1.002462
18499.000000   1.002462
18748.000000   1.002462
18999.000000   1.002462
19249.000000   1.002462
19499.000000   1.002642
19749.000000   1.002642
19999.000000   1.002462
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = No
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 25 October 2019  12:02:56
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 5
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 12:59:55
@@Data
New Section: Section 0: 
2.964000E+1   9.005901E+1   9.005901E+1   9.999000E+3   9.999000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -2.799961E-1   3.513825E-1   -4.019584E-4   -2.263013E-5   2.263013E-5   -4.019584E-4   4.025949E-4   -1.767777E+2   -8.677767E+1   
5.501000E+1   9.001721E+1   9.001721E+1   9.498000E+3   9.498000E+3   9.000000E+1   9.498000E+3   9.498000E+3   -2.481703E-1   3.190423E-1   -3.612193E-4   -2.502638E-5   2.502638E-5   -3.612193E-4   3.620852E-4   -1.760367E+2   -8.603671E+1   
8.006400E+1   9.004751E+1   9.004751E+1   8.998000E+3   8.998000E+3   9.000000E+1   8.998000E+3   8.998000E+3   -2.309322E-1   2.963801E-1   -3.358023E-4   -2.296034E-5   2.296034E-5   -3.358023E-4   3.365863E-4   -1.760885E+2   -8.608851E+1   
1.052510E+2   8.996789E+1   8.996789E+1   8.498000E+3   8.498000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -2.035196E-1   2.666618E-1   -2.994994E-4   -2.380649E-5   2.380649E-5   -2.994994E-4   3.004440E-4   -1.754553E+2   -8.545525E+1   
1.310900E+2   9.003799E+1   9.003799E+1   7.999000E+3   7.999000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -1.790234E-1   2.388935E-1   -2.662694E-4   -2.377054E-5   2.377054E-5   -2.662694E-4   2.673283E-4   -1.748986E+2   -8.489859E+1   
1.568430E+2   8.997659E+1   8.997659E+1   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -1.524067E-1   2.084443E-1   -2.299825E-4   -2.355026E-5   2.355026E-5   -2.299825E-4   2.311851E-4   -1.741533E+2   -8.415328E+1   
1.817480E+2   9.001739E+1   9.001739E+1   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -1.328266E-1   1.824448E-1   -2.009440E-4   -2.103462E-5   2.103462E-5   -2.009440E-4   2.020419E-4   -1.740241E+2   -8.402410E+1   
2.071170E+2   8.993179E+1   8.993179E+1   6.498000E+3   6.498000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -1.126556E-1   1.593506E-1   -1.734323E-4   -2.085537E-5   2.085537E-5   -1.734323E-4   1.746817E-4   -1.731431E+2   -8.314306E+1   
2.325250E+2   8.997680E+1   8.997680E+1   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -9.650652E-2   1.360055E-1   -1.482438E-4   -1.753736E-5   1.753736E-5   -1.482438E-4   1.492776E-4   -1.732532E+2   -8.325322E+1   
2.579260E+2   9.001901E+1   9.001901E+1   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -7.746671E-2   1.137373E-1   -1.219694E-4   -1.706146E-5   1.706146E-5   -1.219694E-4   1.231570E-4   -1.720370E+2   -8.203696E+1   
2.833040E+2   9.000771E+1   9.000771E+1   4.998000E+3   4.998000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -5.860879E-2   8.963229E-2   -9.461126E-5   -1.525018E-5   1.525018E-5   -9.461126E-5   9.583245E-5   -1.708434E+2   -8.084338E+1   
3.084710E+2   9.003619E+1   9.003619E+1   4.497000E+3   4.497000E+3   9.000000E+1   4.498000E+3   4.498000E+3   -4.427347E-2   6.958644E-2   -7.269284E-5   -1.274761E-5   1.274761E-5   -7.269284E-5   7.380211E-5   -1.700536E+2   -8.005359E+1   
3.338730E+2   9.000009E+1   9.000009E+1   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -2.448711E-2   4.660390E-2   -4.549170E-5   -1.235689E-5   1.235689E-5   -4.549170E-5   4.714009E-5   -1.648034E+2   -7.480344E+1   
3.597210E+2   8.997750E+1   8.997750E+1   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -8.998885E-3   2.635550E-2   -2.272859E-5   -1.057463E-5   1.057463E-5   -2.272859E-5   2.506814E-5   -1.550495E+2   -6.504948E+1   
3.847660E+2   9.000411E+1   9.000411E+1   2.998000E+3   2.998000E+3   9.000000E+1   2.998000E+3   2.998000E+3   6.065937E-3   6.171473E-3   -2.691685E-7   -8.521290E-6   8.521290E-6   -2.691685E-7   8.525541E-6   -9.180924E+1   -1.809244E+0   
4.105240E+2   8.999871E+1   8.999871E+1   2.498000E+3   2.498000E+3   9.000000E+1   2.498000E+3   2.498000E+3   2.068039E-2   -1.412911E-2   2.198772E-5   -6.058645E-6   6.058645E-6   2.198772E-5   2.280717E-5   -1.540537E+1   7.459463E+1   
4.363770E+2   9.002801E+1   9.002801E+1   1.998000E+3   1.998000E+3   9.000000E+1   1.999000E+3   1.999000E+3   3.757000E-2   -3.776942E-2   4.782635E-5   -3.095365E-6   3.095365E-6   4.782635E-5   4.792642E-5   -3.703070E+0   8.629693E+1   
4.704600E+2   8.999349E+1   8.999349E+1   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   4.061093E-2   -3.871188E-2   5.032022E-5   -4.728372E-6   4.728372E-6   5.032022E-5   5.054188E-5   -5.368074E+0   8.463193E+1   
4.927400E+2   9.003549E+1   9.003549E+1   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   4.078702E-2   -4.070113E-2   5.172465E-5   -3.558099E-6   3.558099E-6   5.172465E-5   5.184689E-5   -3.935133E+0   8.606487E+1   
5.148310E+2   8.998629E+1   8.998629E+1   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   4.294869E-2   -4.320086E-2   5.468915E-5   -3.522687E-6   3.522687E-6   5.468915E-5   5.480249E-5   -3.685496E+0   8.631450E+1   
5.368250E+2   9.000900E+1   9.000900E+1   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   4.462626E-2   -4.382919E-2   5.613553E-5   -4.352683E-6   4.352683E-6   5.613553E-5   5.630402E-5   -4.433776E+0   8.556622E+1   
5.588170E+2   9.000509E+1   9.000509E+1   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   4.570926E-2   -4.812993E-2   5.960612E-5   -2.342000E-6   2.342000E-6   5.960612E-5   5.965211E-5   -2.250066E+0   8.774993E+1   
5.808840E+2   9.000149E+1   9.000149E+1   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   4.787650E-2   -4.848457E-2   6.117698E-5   -3.713103E-6   3.713103E-6   6.117698E-5   6.128956E-5   -3.473275E+0   8.652673E+1   
6.031090E+2   9.002459E+1   9.002459E+1   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   4.821582E-2   -5.068861E-2   6.282223E-5   -2.523139E-6   2.523139E-6   6.282223E-5   6.287288E-5   -2.299943E+0   8.770006E+1   
6.251690E+2   9.004009E+1   9.004009E+1   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   5.249501E-2   -5.374857E-2   6.746075E-5   -3.687642E-6   3.687642E-6   6.746075E-5   6.756146E-5   -3.128875E+0   8.687113E+1   
6.476280E+2   9.000710E+1   9.000710E+1   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   5.299325E-2   -5.653855E-2   6.958586E-5   -2.232149E-6   2.232149E-6   6.958586E-5   6.962166E-5   -1.837283E+0   8.816272E+1   
6.696560E+2   9.006091E+1   9.006091E+1   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   5.395902E-2   -5.718526E-2   7.060415E-5   -2.523659E-6   2.523659E-6   7.060415E-5   7.064924E-5   -2.047097E+0   8.795290E+1   
6.919480E+2   9.002749E+1   9.002749E+1   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   5.501746E-2   -5.960158E-2   7.283224E-5   -1.726793E-6   1.726793E-6   7.283224E-5   7.285271E-5   -1.358182E+0   8.864182E+1   
7.141830E+2   9.006240E+1   9.006240E+1   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   5.747365E-2   -6.165155E-2   7.568590E-5   -2.203255E-6   2.203255E-6   7.568590E-5   7.571796E-5   -1.667438E+0   8.833256E+1   
7.364830E+2   8.999749E+1   8.999749E+1   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   5.904504E-2   -6.348001E-2   7.784827E-5   -2.170109E-6   2.170109E-6   7.784827E-5   7.787851E-5   -1.596771E+0   8.840323E+1   
7.587120E+2   8.994549E+1   8.994549E+1   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   6.043419E-2   -6.460228E-2   7.943802E-5   -2.463863E-6   2.463863E-6   7.943802E-5   7.947622E-5   -1.776526E+0   8.822347E+1   
7.810190E+2   9.004080E+1   9.004080E+1   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   6.127419E-2   -6.691182E-2   8.146153E-5   -1.575235E-6   1.575235E-6   8.146153E-5   8.147676E-5   -1.107800E+0   8.889220E+1   
8.032580E+2   9.004751E+1   9.004751E+1   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   6.244123E-2   -6.969259E-2   8.399414E-5   -6.204256E-7   6.204256E-7   8.399414E-5   8.399643E-5   -4.232096E-1   8.957679E+1   
8.255590E+2   9.002761E+1   9.002761E+1   1.148000E+3   1.148000E+3   9.000000E+1   1.148000E+3   1.148000E+3   6.293763E-2   -7.065653E-2   8.492883E-5   -3.573814E-7   3.573814E-7   8.492883E-5   8.492959E-5   -2.410998E-1   8.975890E+1   
8.479080E+2   9.008209E+1   9.008209E+1   1.097000E+3   1.097000E+3   9.000000E+1   1.098000E+3   1.098000E+3   6.543430E-2   -7.298508E-2   8.798895E-5   -6.816564E-7   6.816564E-7   8.798895E-5   8.799159E-5   -4.438654E-1   8.955613E+1   
8.701470E+2   9.005190E+1   9.005190E+1   1.047000E+3   1.047000E+3   9.000000E+1   1.048000E+3   1.048000E+3   6.664184E-2   -7.546581E-2   9.035119E-5   4.704014E-8   -4.704014E-8   9.035119E-5   9.035120E-5   2.983028E-2   9.002983E+1   
8.922800E+2   9.000079E+1   9.000079E+1   9.980000E+2   9.980000E+2   9.000000E+1   9.990000E+2   9.990000E+2   7.014665E-2   -7.729921E-2   9.371209E-5   -1.346604E-6   1.346604E-6   9.371209E-5   9.372177E-5   -8.232597E-1   8.917674E+1   
9.142010E+2   9.000521E+1   9.000521E+1   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   7.104616E-2   -7.973145E-2   9.585231E-5   -4.217772E-7   4.217772E-7   9.585231E-5   9.585324E-5   -2.521160E-1   8.974788E+1   
9.360780E+2   9.000720E+1   9.000720E+1   8.980000E+2   8.980000E+2   9.000000E+1   8.980000E+2   8.980000E+2   7.186651E-2   -8.184587E-2   9.773658E-5   3.538133E-7   -3.538133E-7   9.773658E-5   9.773722E-5   2.074139E-1   9.020741E+1   
9.579550E+2   9.001739E+1   9.001739E+1   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   7.276788E-2   -8.429777E-2   9.989075E-5   1.290116E-6   -1.290116E-6   9.989075E-5   9.989908E-5   7.399495E-1   9.073995E+1   
9.798280E+2   9.007250E+1   9.007250E+1   7.980000E+2   7.980000E+2   9.000000E+1   7.990000E+2   7.990000E+2   7.612481E-2   -8.605626E-2   1.031114E-4   -4.311929E-8   4.311929E-8   1.031114E-4   1.031115E-4   -2.396003E-2   8.997604E+1   
1.001696E+3   8.999691E+1   8.999691E+1   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   7.773913E-2   -8.755405E-2   1.050850E-4   -2.579153E-7   2.579153E-7   1.050850E-4   1.050853E-4   -1.406236E-1   8.985938E+1   
1.023543E+3   9.000329E+1   9.000329E+1   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   7.905039E-2   -8.908250E-2   1.068911E-4   -2.285037E-7   2.285037E-7   1.068911E-4   1.068914E-4   -1.224824E-1   8.987752E+1   
1.045439E+3   8.997659E+1   8.997659E+1   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   8.049658E-2   -9.087907E-2   1.089553E-4   -1.236067E-7   1.236067E-7   1.089553E-4   1.089554E-4   -6.500037E-2   8.993500E+1   
1.067310E+3   8.999291E+1   8.999291E+1   5.980000E+2   5.980000E+2   9.000000E+1   5.990000E+2   5.990000E+2   8.040210E-2   -9.264995E-2   1.100503E-4   1.104023E-6   -1.104023E-6   1.100503E-4   1.100558E-4   5.747716E-1   9.057477E+1   
1.089177E+3   8.999490E+1   8.999490E+1   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   8.055611E-2   -9.477247E-2   1.115279E-4   2.377762E-6   -2.377762E-6   1.115279E-4   1.115532E-4   1.221355E+0   9.122135E+1   
1.111000E+3   9.002761E+1   9.002761E+1   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   8.311967E-2   -9.696491E-2   1.145407E-4   1.915029E-6   -1.915029E-6   1.145407E-4   1.145567E-4   9.578504E-1   9.095785E+1   
1.132896E+3   9.002340E+1   9.002340E+1   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   8.534145E-2   -9.871488E-2   1.170540E-4   1.415810E-6   -1.415810E-6   1.170540E-4   1.170626E-4   6.929789E-1   9.069298E+1   
1.154778E+3   9.001211E+1   9.001211E+1   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   8.463094E-2   -1.003722E-1   1.176942E-4   3.024840E-6   -3.024840E-6   1.176942E-4   1.177330E-4   1.472226E+0   9.147223E+1   
1.176666E+3   8.996270E+1   8.996270E+1   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   8.667784E-2   -1.026694E-1   1.204558E-4   3.012763E-6   -3.012763E-6   1.204558E-4   1.204935E-4   1.432746E+0   9.143275E+1   
1.198491E+3   9.000720E+1   9.000720E+1   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   8.936104E-2   -1.047912E-1   1.234966E-4   2.415357E-6   -2.415357E-6   1.234966E-4   1.235202E-4   1.120453E+0   9.112045E+1   
1.220328E+3   9.001809E+1   9.001809E+1   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   8.935921E-2   -1.061049E-1   1.243511E-4   3.275548E-6   -3.275548E-6   1.243511E-4   1.243942E-4   1.508887E+0   9.150889E+1   
1.242097E+3   9.003259E+1   9.003259E+1   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   9.165836E-2   -1.071413E-1   1.264475E-4   2.252571E-6   -2.252571E-6   1.264475E-4   1.264675E-4   1.020575E+0   9.102058E+1   
1.263929E+3   9.003561E+1   9.003561E+1   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   9.342864E-2   -1.103098E-1   1.296056E-4   3.014733E-6   -3.014733E-6   1.296056E-4   1.296406E-4   1.332507E+0   9.133251E+1   
1.285748E+3   9.005139E+1   9.005139E+1   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   9.433192E-2   -1.113885E-1   1.308666E-4   3.051835E-6   -3.051835E-6   1.308666E-4   1.309021E-4   1.335907E+0   9.133591E+1   
1.307477E+3   9.004681E+1   9.004681E+1   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   9.409014E-2   -1.143834E-1   1.326676E-4   5.188657E-6   -5.188657E-6   1.326676E-4   1.327691E-4   2.239708E+0   9.223971E+1   
1.340666E+3   9.003039E+1   9.003039E+1   4.600000E+1   4.600000E+1   9.000000E+1   4.700000E+1   4.700000E+1   9.547567E-2   -1.139306E-1   1.332293E-4   3.867831E-6   -3.867831E-6   1.332293E-4   1.332854E-4   1.662909E+0   9.166291E+1   
1.359747E+3   9.000610E+1   9.000610E+1   4.600000E+1   4.600000E+1   9.000000E+1   4.700000E+1   4.700000E+1   9.564623E-2   -1.134937E-1   1.330502E-4   3.456069E-6   -3.456069E-6   1.330502E-4   1.330951E-4   1.487962E+0   9.148796E+1   
1.382177E+3   9.002831E+1   9.002831E+1   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   9.564627E-2   -1.134784E-1   1.330403E-4   3.445995E-6   -3.445995E-6   1.330403E-4   1.330849E-4   1.483737E+0   9.148374E+1   
1.401281E+3   8.999841E+1   8.999841E+1   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   9.586536E-2   -1.132084E-1   1.329999E-4   3.107452E-6   -3.107452E-6   1.329999E-4   1.330362E-4   1.338434E+0   9.133843E+1   
1.423687E+3   9.000771E+1   9.000771E+1   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   9.612796E-2   -1.127439E-1   1.328597E-4   2.609556E-6   -2.609556E-6   1.328597E-4   1.328853E-4   1.125227E+0   9.112523E+1   
1.442739E+3   8.999240E+1   8.999240E+1   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   9.540142E-2   -1.127003E-1   1.323822E-4   3.118451E-6   -3.118451E-6   1.323822E-4   1.324189E-4   1.349434E+0   9.134943E+1   
1.465105E+3   9.001870E+1   9.001870E+1   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   9.545361E-2   -1.144319E-1   1.335422E-4   4.211877E-6   -4.211877E-6   1.335422E-4   1.336086E-4   1.806491E+0   9.180649E+1   
1.484178E+3   9.002221E+1   9.002221E+1   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   9.617272E-2   -1.141772E-1   1.338209E-4   3.513528E-6   -3.513528E-6   1.338209E-4   1.338670E-4   1.503981E+0   9.150398E+1   
1.506619E+3   8.998821E+1   8.998821E+1   3.000000E+1   3.000000E+1   9.000000E+1   3.100000E+1   3.100000E+1   9.751714E-2   -1.138570E-1   1.344435E-4   2.309763E-6   -2.309763E-6   1.344435E-4   1.344633E-4   9.842548E-1   9.098425E+1   
1.525712E+3   9.002331E+1   9.002331E+1   3.000000E+1   3.000000E+1   9.000000E+1   3.100000E+1   3.100000E+1   9.665379E-2   -1.142012E-1   1.341339E-4   3.173356E-6   -3.173356E-6   1.341339E-4   1.341714E-4   1.355257E+0   9.135526E+1   
1.548134E+3   9.002291E+1   9.002291E+1   2.600000E+1   2.600000E+1   9.000000E+1   2.700000E+1   2.700000E+1   9.593037E-2   -1.147080E-1   1.340167E-4   4.039767E-6   -4.039767E-6   1.340167E-4   1.340776E-4   1.726587E+0   9.172659E+1   
1.567162E+3   9.002981E+1   9.002981E+1   2.600000E+1   2.600000E+1   9.000000E+1   2.700000E+1   2.700000E+1   9.557389E-2   -1.137202E-1   1.331530E-4   3.657603E-6   -3.657603E-6   1.331530E-4   1.332032E-4   1.573472E+0   9.157347E+1   
1.589589E+3   9.003091E+1   9.003091E+1   2.200000E+1   2.200000E+1   9.000000E+1   2.300000E+1   2.300000E+1   9.647221E-2   -1.138852E-1   1.338158E-4   3.101066E-6   -3.101066E-6   1.338158E-4   1.338518E-4   1.327542E+0   9.132754E+1   
1.608677E+3   8.996691E+1   8.996691E+1   2.200000E+1   2.200000E+1   9.000000E+1   2.300000E+1   2.300000E+1   9.582851E-2   -1.136913E-1   1.332916E-4   3.450402E-6   -3.450402E-6   1.332916E-4   1.333362E-4   1.482834E+0   9.148283E+1   
1.631072E+3   9.000689E+1   9.000689E+1   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   9.659242E-2   -1.147141E-1   1.344301E-4   3.554110E-6   -3.554110E-6   1.344301E-4   1.344770E-4   1.514454E+0   9.151445E+1   
1.650063E+3   9.005389E+1   9.005389E+1   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   9.768592E-2   -1.147086E-1   1.351025E-4   2.741710E-6   -2.741710E-6   1.351025E-4   1.351303E-4   1.162576E+0   9.116258E+1   
1.672453E+3   9.002349E+1   9.002349E+1   1.500000E+1   1.500000E+1   9.000000E+1   1.500000E+1   1.500000E+1   9.656301E-2   -1.141239E-1   1.340274E-4   3.189959E-6   -3.189959E-6   1.340274E-4   1.340654E-4   1.363428E+0   9.136343E+1   
1.693876E+3   9.002542E+1   9.002542E+1   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   9.684708E-2   -1.150620E-1   1.348141E-4   3.593202E-6   -3.593202E-6   1.348141E-4   1.348620E-4   1.526744E+0   9.152674E+1   
1.712953E+3   8.997341E+1   8.997341E+1   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   9.610035E-2   -1.142318E-1   1.338117E-4   3.602747E-6   -3.602747E-6   1.338117E-4   1.338602E-4   1.542259E+0   9.154226E+1   
1.735079E+3   9.001650E+1   9.001650E+1   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   9.530876E-2   -1.145804E-1   1.335493E-4   4.416097E-6   -4.416097E-6   1.335493E-4   1.336223E-4   1.893919E+0   9.189392E+1   
1.753792E+3   9.003030E+1   9.003030E+1   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   9.788527E-2   -1.151424E-1   1.355083E-4   2.877874E-6   -2.877874E-6   1.355083E-4   1.355388E-4   1.216643E+0   9.121664E+1   
1.775791E+3   8.998940E+1   8.998940E+1   5.000000E+0   5.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   9.711892E-2   -1.145976E-1   1.346796E-4   3.088472E-6   -3.088472E-6   1.346796E-4   1.347150E-4   1.313676E+0   9.131368E+1   
1.796771E+3   9.001989E+1   9.001989E+1   3.000000E+0   3.000000E+0   9.000000E+1   3.000000E+0   3.000000E+0   9.690660E-2   -1.147006E-1   1.346155E-4   3.312907E-6   -3.312907E-6   1.346155E-4   1.346563E-4   1.409773E+0   9.140977E+1   
1.817854E+3   9.005050E+1   9.005050E+1   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   9.637460E-2   -1.145681E-1   1.342003E-4   3.619750E-6   -3.619750E-6   1.342003E-4   1.342491E-4   1.545050E+0   9.154505E+1   
1.836571E+3   9.000939E+1   9.000939E+1   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   9.653170E-2   -1.153836E-1   1.348285E-4   4.036685E-6   -4.036685E-6   1.348285E-4   1.348889E-4   1.714889E+0   9.171489E+1   
1.858572E+3   9.006951E+1   9.006951E+1   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   9.676304E-2   -1.160002E-1   1.353731E-4   4.268705E-6   -4.268705E-6   1.353731E-4   1.354404E-4   1.806103E+0   9.180610E+1   
1.880613E+3   9.000701E+1   9.000701E+1   -3.000000E+0   -3.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   9.729566E-2   -1.161420E-1   1.357948E-4   3.967434E-6   -3.967434E-6   1.357948E-4   1.358527E-4   1.673501E+0   9.167350E+1   
1.902404E+3   9.001559E+1   9.001559E+1   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   9.697532E-2   -1.146951E-1   1.346544E-4   3.258458E-6   -3.258458E-6   1.346544E-4   1.346938E-4   1.386212E+0   9.138621E+1   
1.924471E+3   9.004379E+1   9.004379E+1   -8.000000E+0   -8.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   9.703979E-2   -1.158284E-1   1.354324E-4   3.951706E-6   -3.951706E-6   1.354324E-4   1.354900E-4   1.671328E+0   9.167133E+1   
1.946523E+3   9.000689E+1   9.000689E+1   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   9.726619E-2   -1.158057E-1   1.355575E-4   3.769406E-6   -3.769406E-6   1.355575E-4   1.356099E-4   1.592795E+0   9.159280E+1   
1.968793E+3   9.003460E+1   9.003460E+1   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   9.748893E-2   -1.156100E-1   1.355678E-4   3.476691E-6   -3.476691E-6   1.355678E-4   1.356123E-4   1.469052E+0   9.146905E+1   
1.991002E+3   9.005929E+1   9.005929E+1   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   9.696371E-2   -1.154639E-1   1.351479E-4   3.769690E-6   -3.769690E-6   1.351479E-4   1.352005E-4   1.597741E+0   9.159774E+1   
2.013233E+3   9.003771E+1   9.003771E+1   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   9.803258E-2   -1.160947E-1   1.362196E-4   3.391494E-6   -3.391494E-6   1.362196E-4   1.362618E-4   1.426213E+0   9.142621E+1   
2.035507E+3   8.999731E+1   8.999731E+1   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   9.681152E-2   -1.167396E-1   1.358847E-4   4.716224E-6   -4.716224E-6   1.358847E-4   1.359665E-4   1.987798E+0   9.198780E+1   
2.057754E+3   8.995791E+1   8.995791E+1   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   9.801353E-2   -1.162383E-1   1.363013E-4   3.499449E-6   -3.499449E-6   1.363013E-4   1.363462E-4   1.470710E+0   9.147071E+1   
2.079995E+3   8.996761E+1   8.996761E+1   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   9.781844E-2   -1.163223E-1   1.362354E-4   3.698694E-6   -3.698694E-6   1.362354E-4   1.362856E-4   1.555157E+0   9.155516E+1   
2.102217E+3   9.002221E+1   9.002221E+1   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   9.783257E-2   -1.168997E-1   1.366202E-4   4.065732E-6   -4.065732E-6   1.366202E-4   1.366807E-4   1.704583E+0   9.170458E+1   
2.124456E+3   8.998699E+1   8.998699E+1   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   9.734902E-2   -1.164359E-1   1.360192E-4   4.120122E-6   -4.120122E-6   1.360192E-4   1.360815E-4   1.735002E+0   9.173500E+1   
2.146637E+3   9.000079E+1   9.000079E+1   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   9.718579E-2   -1.159708E-1   1.356153E-4   3.936778E-6   -3.936778E-6   1.356153E-4   1.356725E-4   1.662772E+0   9.166277E+1   
2.168910E+3   9.000469E+1   9.000469E+1   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   9.767670E-2   -1.159198E-1   1.358857E-4   3.540387E-6   -3.540387E-6   1.358857E-4   1.359318E-4   1.492456E+0   9.149246E+1   
2.191181E+3   8.996899E+1   8.996899E+1   -3.100000E+1   -3.100000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   9.794973E-2   -1.162886E-1   1.362946E-4   3.579534E-6   -3.579534E-6   1.362946E-4   1.363416E-4   1.504425E+0   9.150442E+1   
2.213132E+3   9.003671E+1   9.003671E+1   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   9.706247E-2   -1.175133E-1   1.365437E-4   5.036467E-6   -5.036467E-6   1.365437E-4   1.366366E-4   2.112419E+0   9.211242E+1   
2.235370E+3   8.996179E+1   8.996179E+1   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   9.941685E-2   -1.161800E-1   1.371309E-4   2.423416E-6   -2.423416E-6   1.371309E-4   1.371524E-4   1.012442E+0   9.101244E+1   
2.257611E+3   9.002859E+1   9.002859E+1   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   9.748404E-2   -1.171838E-1   1.365898E-4   4.509249E-6   -4.509249E-6   1.365898E-4   1.366642E-4   1.890823E+0   9.189082E+1   
2.279855E+3   9.000390E+1   9.000390E+1   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   9.830134E-2   -1.164322E-1   1.366055E-4   3.413336E-6   -3.413336E-6   1.366055E-4   1.366482E-4   1.431341E+0   9.143134E+1   
2.302117E+3   9.006671E+1   9.006671E+1   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   9.747790E-2   -1.172777E-1   1.366471E-4   4.575160E-6   -4.575160E-6   1.366471E-4   1.367237E-4   1.917636E+0   9.191764E+1   
2.324400E+3   9.003741E+1   9.003741E+1   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   9.726251E-2   -1.174826E-1   1.366474E-4   4.868460E-6   -4.868460E-6   1.366474E-4   1.367341E-4   2.040465E+0   9.204046E+1   
2.346678E+3   8.997189E+1   8.997189E+1   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   9.794053E-2   -1.168758E-1   1.366714E-4   3.970236E-6   -3.970236E-6   1.366714E-4   1.367290E-4   1.663946E+0   9.166395E+1   
2.368951E+3   9.002551E+1   9.002551E+1   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   9.923031E-2   -1.170758E-1   1.375991E-4   3.147056E-6   -3.147056E-6   1.375991E-4   1.376351E-4   1.310195E+0   9.131019E+1   
2.391210E+3   8.999749E+1   8.999749E+1   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   9.787428E-2   -1.177692E-1   1.372123E-4   4.603296E-6   -4.603296E-6   1.372123E-4   1.372895E-4   1.921479E+0   9.192148E+1   
2.424527E+3   9.007479E+1   9.007479E+1   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   9.978745E-2   -1.187215E-1   1.390153E-4   3.810845E-6   -3.810845E-6   1.390153E-4   1.390675E-4   1.570264E+0   9.157026E+1   
2.446268E+3   9.001650E+1   9.001650E+1   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   1.014779E-1   -1.202223E-1   1.410379E-4   3.541765E-6   -3.541765E-6   1.410379E-4   1.410823E-4   1.438518E+0   9.143852E+1   
2.467984E+3   9.003701E+1   9.003701E+1   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   1.022786E-1   -1.226834E-1   1.431358E-4   4.558478E-6   -4.558478E-6   1.431358E-4   1.432084E-4   1.824095E+0   9.182409E+1   
2.489679E+3   9.001199E+1   9.001199E+1   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   1.028768E-1   -1.239934E-1   1.443589E-4   4.972465E-6   -4.972465E-6   1.443589E-4   1.444445E-4   1.972783E+0   9.197278E+1   
2.511844E+3   9.000509E+1   9.000509E+1   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   1.059037E-1   -1.259372E-1   1.474962E-4   4.004549E-6   -4.004549E-6   1.474962E-4   1.475505E-4   1.555209E+0   9.155521E+1   
2.533513E+3   8.996200E+1   8.996200E+1   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   1.074751E-1   -1.283535E-1   1.500414E-4   4.422019E-6   -4.422019E-6   1.500414E-4   1.501065E-4   1.688132E+0   9.168813E+1   
2.555232E+3   9.002490E+1   9.002490E+1   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   1.088753E-1   -1.289763E-1   1.513127E-4   3.793550E-6   -3.793550E-6   1.513127E-4   1.513602E-4   1.436158E+0   9.143616E+1   
2.577607E+3   9.001989E+1   9.001989E+1   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   1.086188E-1   -1.309570E-1   1.524441E-4   5.278134E-6   -5.278134E-6   1.524441E-4   1.525354E-4   1.982983E+0   9.198298E+1   
2.599256E+3   9.002499E+1   9.002499E+1   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   1.091195E-1   -1.327235E-1   1.539042E-4   6.062714E-6   -6.062714E-6   1.539042E-4   1.540235E-4   2.255874E+0   9.225587E+1   
2.620928E+3   9.000179E+1   9.000179E+1   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   1.117211E-1   -1.334555E-1   1.559893E-4   4.617057E-6   -4.617057E-6   1.559893E-4   1.560577E-4   1.695377E+0   9.169538E+1   
2.642618E+3   9.002490E+1   9.002490E+1   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   1.139153E-1   -1.363412E-1   1.592253E-4   4.880742E-6   -4.880742E-6   1.592253E-4   1.593001E-4   1.755741E+0   9.175574E+1   
2.664329E+3   8.998190E+1   8.998190E+1   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.500000E+2   -6.500000E+2   1.141306E-1   -1.375407E-1   1.601397E-4   5.505700E-6   -5.505700E-6   1.601397E-4   1.602343E-4   1.969088E+0   9.196909E+1   
2.686008E+3   9.008499E+1   9.008499E+1   -7.010000E+2   -7.010000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   1.153559E-1   -1.395263E-1   1.621904E-4   5.897533E-6   -5.897533E-6   1.621904E-4   1.622976E-4   2.082459E+0   9.208246E+1   
2.707698E+3   8.997521E+1   8.997521E+1   -7.510000E+2   -7.510000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   1.157940E-1   -1.416947E-1   1.638736E-4   6.991120E-6   -6.991120E-6   1.638736E-4   1.640226E-4   2.442852E+0   9.244285E+1   
2.729417E+3   9.000390E+1   9.000390E+1   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   1.173881E-1   -1.430495E-1   1.657415E-4   6.697815E-6   -6.697815E-6   1.657415E-4   1.658768E-4   2.314133E+0   9.231413E+1   
2.751111E+3   9.001879E+1   9.001879E+1   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   1.185926E-1   -1.438085E-1   1.669805E-4   6.303148E-6   -6.303148E-6   1.669805E-4   1.670994E-4   2.161764E+0   9.216176E+1   
2.772840E+3   9.000570E+1   9.000570E+1   -9.000000E+2   -9.000000E+2   9.000000E+1   -8.990000E+2   -8.990000E+2   1.194418E-1   -1.457818E-1   1.687907E-4   6.965162E-6   -6.965162E-6   1.687907E-4   1.689343E-4   2.362975E+0   9.236297E+1   
2.794539E+3   8.999340E+1   8.999340E+1   -9.510000E+2   -9.510000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   1.200585E-1   -1.487423E-1   1.711001E-4   8.444565E-6   -8.444565E-6   1.711001E-4   1.713083E-4   2.825514E+0   9.282551E+1   
2.816226E+3   8.997219E+1   8.997219E+1   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   1.215863E-1   -1.489921E-1   1.722073E-4   7.477820E-6   -7.477820E-6   1.722073E-4   1.723696E-4   2.486414E+0   9.248641E+1   
2.838294E+3   9.005190E+1   9.005190E+1   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   1.238338E-1   -1.504033E-1   1.745160E-4   6.738084E-6   -6.738084E-6   1.745160E-4   1.746460E-4   2.211099E+0   9.221110E+1   
2.860081E+3   9.003860E+1   9.003860E+1   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   1.241333E-1   -1.536713E-1   1.768295E-4   8.653107E-6   -8.653107E-6   1.768295E-4   1.770411E-4   2.801520E+0   9.280152E+1   
2.881923E+3   9.001830E+1   9.001830E+1   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   1.249064E-1   -1.542345E-1   1.776743E-4   8.449530E-6   -8.449530E-6   1.776743E-4   1.778751E-4   2.722723E+0   9.272272E+1   
2.904565E+3   9.001251E+1   9.001251E+1   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   1.262201E-1   -1.564269E-1   1.799143E-4   8.911182E-6   -8.911182E-6   1.799143E-4   1.801349E-4   2.835551E+0   9.283555E+1   
2.926605E+3   9.001281E+1   9.001281E+1   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   1.283247E-1   -1.579565E-1   1.822117E-4   8.354610E-6   -8.354610E-6   1.822117E-4   1.824032E-4   2.625236E+0   9.262524E+1   
2.948734E+3   8.998751E+1   8.998751E+1   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   1.297065E-1   -1.604698E-1   1.847029E-4   8.975684E-6   -8.975684E-6   1.847029E-4   1.849208E-4   2.782115E+0   9.278211E+1   
2.971080E+3   9.008929E+1   9.008929E+1   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   1.308570E-1   -1.610877E-1   1.858166E-4   8.528696E-6   -8.528696E-6   1.858166E-4   1.860122E-4   2.627944E+0   9.262794E+1   
2.993148E+3   9.006429E+1   9.006429E+1   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   1.319240E-1   -1.635770E-1   1.880975E-4   9.366941E-6   -9.366941E-6   1.880975E-4   1.883306E-4   2.850879E+0   9.285088E+1   
3.015269E+3   9.006921E+1   9.006921E+1   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   1.333278E-1   -1.671861E-1   1.913160E-4   1.068813E-5   -1.068813E-5   1.913160E-4   1.916143E-4   3.197583E+0   9.319758E+1   
3.037623E+3   9.001730E+1   9.001730E+1   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   1.344568E-1   -1.678752E-1   1.924628E-4   1.030358E-5   -1.030358E-5   1.924628E-4   1.927384E-4   3.064428E+0   9.306443E+1   
3.059664E+3   9.005770E+1   9.005770E+1   -1.550000E+3   -1.550000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   1.350956E-1   -1.692404E-1   1.937469E-4   1.072369E-5   -1.072369E-5   1.937469E-4   1.940434E-4   3.168029E+0   9.316803E+1   
3.081791E+3   8.999441E+1   8.999441E+1   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   1.360454E-1   -1.712370E-1   1.956345E-4   1.132649E-5   -1.132649E-5   1.956345E-4   1.959621E-4   3.313508E+0   9.331351E+1   
3.104666E+3   9.001599E+1   9.001599E+1   -1.650000E+3   -1.650000E+3   9.000000E+1   -1.648000E+3   -1.648000E+3   1.377450E-1   -1.727955E-1   1.977003E-4   1.108831E-5   -1.108831E-5   1.977003E-4   1.980110E-4   3.210153E+0   9.321015E+1   
3.126739E+3   9.002831E+1   9.002831E+1   -1.700000E+3   -1.700000E+3   9.000000E+1   -1.698000E+3   -1.698000E+3   1.394680E-1   -1.757321E-1   2.006781E-4   1.173384E-5   -1.173384E-5   2.006781E-4   2.010208E-4   3.346328E+0   9.334633E+1   
3.148880E+3   8.999850E+1   8.999850E+1   -1.750000E+3   -1.750000E+3   9.000000E+1   -1.748000E+3   -1.748000E+3   1.397239E-1   -1.773139E-1   2.018665E-4   1.257874E-5   -1.257874E-5   2.018665E-4   2.022580E-4   3.565613E+0   9.356561E+1   
3.171715E+3   9.002490E+1   9.002490E+1   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.798000E+3   -1.798000E+3   1.405516E-1   -1.775729E-1   2.025469E-4   1.213579E-5   -1.213579E-5   2.025469E-4   2.029101E-4   3.428833E+0   9.342883E+1   
3.193819E+3   9.000521E+1   9.000521E+1   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.848000E+3   -1.848000E+3   1.438367E-1   -1.791854E-1   2.056281E-4   1.076023E-5   -1.076023E-5   2.056281E-4   2.059095E-4   2.995475E+0   9.299548E+1   
3.215990E+3   8.999600E+1   8.999600E+1   -1.900000E+3   -1.900000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   1.435674E-1   -1.806954E-1   2.064451E-4   1.194667E-5   -1.194667E-5   2.064451E-4   2.067904E-4   3.311928E+0   9.331193E+1   
3.238828E+3   8.998440E+1   8.998440E+1   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   1.447639E-1   -1.829055E-1   2.086242E-4   1.250663E-5   -1.250663E-5   2.086242E-4   2.089988E-4   3.430667E+0   9.343067E+1   
3.261361E+3   9.008080E+1   9.008080E+1   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   1.471446E-1   -1.844843E-1   2.111243E-4   1.177795E-5   -1.177795E-5   2.111243E-4   2.114526E-4   3.193038E+0   9.319304E+1   
3.298372E+3   9.006289E+1   9.006289E+1   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.594408E-1   -2.037368E-1   2.312654E-4   1.527000E-5   -1.527000E-5   2.312654E-4   2.317690E-4   3.777645E+0   9.377765E+1   
3.324829E+3   9.005190E+1   9.005190E+1   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.720371E-1   -2.228887E-1   2.515264E-4   1.847435E-5   -1.847435E-5   2.515264E-4   2.522040E-4   4.200772E+0   9.420077E+1   
3.349971E+3   9.004199E+1   9.004199E+1   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.853588E-1   -2.422768E-1   2.723897E-4   2.129660E-5   -2.129660E-5   2.723897E-4   2.732210E-4   4.470537E+0   9.447054E+1   
3.375621E+3   8.997451E+1   8.997451E+1   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   1.991319E-1   -2.609082E-1   2.930394E-4   2.329029E-5   -2.329029E-5   2.930394E-4   2.939635E-4   4.544221E+0   9.454422E+1   
3.401776E+3   9.003951E+1   9.003951E+1   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   2.083393E-1   -2.760044E-1   3.085638E-4   2.634961E-5   -2.634961E-5   3.085638E-4   3.096868E-4   4.880894E+0   9.488089E+1   
3.427020E+3   9.000759E+1   9.000759E+1   -5.000000E+3   -5.000000E+3   9.000000E+1   -5.000000E+3   -5.000000E+3   2.138647E-1   -2.844404E-1   3.174742E-4   2.777812E-5   -2.777812E-5   3.174742E-4   3.186871E-4   5.000489E+0   9.500049E+1   
3.452189E+3   9.002590E+1   9.002590E+1   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   2.099132E-1   -2.811461E-1   3.128856E-4   2.854705E-5   -2.854705E-5   3.128856E-4   3.141852E-4   5.213118E+0   9.521312E+1   
3.478360E+3   9.003961E+1   9.003961E+1   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   1.979152E-1   -2.715282E-1   2.992038E-4   3.113323E-5   -3.113323E-5   2.992038E-4   3.008192E-4   5.940454E+0   9.594045E+1   
3.503035E+3   8.997729E+1   8.997729E+1   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.865836E-1   -2.559678E-1   2.820638E-4   2.934151E-5   -2.934151E-5   2.820638E-4   2.835858E-4   5.938798E+0   9.593880E+1   
3.527719E+3   9.001019E+1   9.001019E+1   -7.000000E+3   -7.000000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.775612E-1   -2.453293E-1   2.695570E-4   2.905956E-5   -2.905956E-5   2.695570E-4   2.711189E-4   6.153002E+0   9.615300E+1   
3.552408E+3   9.006451E+1   9.006451E+1   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.729618E-1   -2.408189E-1   2.637759E-4   2.951269E-5   -2.951269E-5   2.637759E-4   2.654217E-4   6.384015E+0   9.638401E+1   
3.578014E+3   9.003469E+1   9.003469E+1   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.999000E+3   -7.999000E+3   1.789608E-1   -2.476881E-1   2.719585E-4   2.956650E-5   -2.956650E-5   2.719585E-4   2.735610E-4   6.204653E+0   9.620465E+1   
3.603265E+3   9.001150E+1   9.001150E+1   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.812115E-1   -2.563273E-1   2.789767E-4   3.354992E-5   -3.354992E-5   2.789767E-4   2.809868E-4   6.857497E+0   9.685750E+1   
3.628950E+3   8.998229E+1   8.998229E+1   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.943513E-1   -2.709889E-1   2.966493E-4   3.341662E-5   -3.341662E-5   2.966493E-4   2.985255E-4   6.427097E+0   9.642710E+1   
3.654143E+3   8.996789E+1   8.996789E+1   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   2.083608E-1   -2.897350E-1   3.175197E-4   3.531040E-5   -3.531040E-5   3.175197E-4   3.194771E-4   6.345615E+0   9.634562E+1   
3.679334E+3   9.002429E+1   9.002429E+1   -9.999000E+3   -9.999000E+3   9.000000E+1   -9.999000E+3   -9.999000E+3   2.178923E-1   -3.066185E-1   3.344086E-4   3.929863E-5   -3.929863E-5   3.344086E-4   3.367098E-4   6.702476E+0   9.670248E+1   
3.715438E+3   9.007940E+1   9.007940E+1   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.956356E-1   -2.761386E-1   3.007972E-4   3.583344E-5   -3.583344E-5   3.007972E-4   3.029241E-4   6.793528E+0   9.679353E+1   
3.739670E+3   9.002679E+1   9.002679E+1   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.717088E-1   -2.496072E-1   2.687250E-4   3.618494E-5   -3.618494E-5   2.687250E-4   2.711502E-4   7.668987E+0   9.766899E+1   
3.764420E+3   9.003130E+1   9.003130E+1   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.568042E-1   -2.298516E-1   2.466436E-4   3.429323E-5   -3.429323E-5   2.466436E-4   2.490163E-4   7.915633E+0   9.791563E+1   
3.789069E+3   9.003979E+1   9.003979E+1   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.434999E-1   -2.122823E-1   2.269755E-4   3.264718E-5   -3.264718E-5   2.269755E-4   2.293114E-4   8.185039E+0   9.818504E+1   
3.813813E+3   8.997109E+1   8.997109E+1   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.279265E-1   -1.905936E-1   2.032217E-4   2.998636E-5   -2.998636E-5   2.032217E-4   2.054221E-4   8.393703E+0   9.839370E+1   
3.839004E+3   9.000219E+1   9.000219E+1   -7.000000E+3   -7.000000E+3   9.000000E+1   -6.999000E+3   -6.999000E+3   1.157266E-1   -1.727801E-1   1.840775E-4   2.736382E-5   -2.736382E-5   1.840775E-4   1.861002E-4   8.455318E+0   9.845532E+1   
3.863741E+3   9.001760E+1   9.001760E+1   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.003973E-1   -1.528711E-1   1.616337E-4   2.568584E-5   -2.568584E-5   1.616337E-4   1.636619E-4   9.029592E+0   9.902959E+1   
3.887993E+3   9.001571E+1   9.001571E+1   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   8.493833E-2   -1.307490E-1   1.376683E-4   2.265694E-5   -2.265694E-5   1.376683E-4   1.395202E-4   9.345755E+0   9.934575E+1   
3.912632E+3   9.003240E+1   9.003240E+1   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   7.295686E-2   -1.135311E-1   1.190470E-4   2.026230E-5   -2.026230E-5   1.190470E-4   1.207590E-4   9.659417E+0   9.965942E+1   
3.937316E+3   9.000100E+1   9.000100E+1   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   5.754666E-2   -9.358878E-2   9.653142E-5   1.862240E-5   -1.862240E-5   9.653142E-5   9.831128E-5   1.091910E+1   1.009191E+2   
3.961530E+3   9.001110E+1   9.001110E+1   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   4.594488E-2   -7.576830E-2   7.775236E-5   1.555291E-5   -1.555291E-5   7.775236E-5   7.929264E-5   1.131166E+1   1.013117E+2   
3.986233E+3   9.005621E+1   9.005621E+1   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   3.452540E-2   -5.704967E-2   5.850106E-5   1.176141E-5   -1.176141E-5   5.850106E-5   5.967164E-5   1.136755E+1   1.013675E+2   
4.010921E+3   9.000930E+1   9.000930E+1   -3.499000E+3   -3.499000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.905130E-2   -3.783016E-2   3.641679E-5   1.064135E-5   -1.064135E-5   3.641679E-5   3.793970E-5   1.628890E+1   1.062889E+2   
4.035594E+3   9.005261E+1   9.005261E+1   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   6.980183E-3   -2.180079E-2   1.851410E-5   9.089983E-6   -9.089983E-6   1.851410E-5   2.062522E-5   2.614994E+1   1.161499E+2   
4.060227E+3   8.999551E+1   8.999551E+1   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   -6.829856E-3   -1.541948E-3   -3.218282E-6   6.059656E-6   -6.059656E-6   -3.218282E-6   6.861251E-6   1.179728E+2   2.079728E+2   
4.084912E+3   9.006680E+1   9.006680E+1   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   -1.976185E-2   1.805238E-2   -2.397502E-5   2.814339E-6   -2.814339E-6   -2.397502E-5   2.413964E-5   1.733049E+2   2.633049E+2   
4.118578E+3   9.003759E+1   9.003759E+1   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   -2.034720E-2   2.212048E-2   -2.698642E-5   5.876767E-7   -5.876767E-7   -2.698642E-5   2.699282E-5   1.787525E+2   2.687525E+2   
4.140608E+3   9.004711E+1   9.004711E+1   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.899000E+3   -1.899000E+3   -2.212293E-2   2.331452E-2   -2.886193E-5   1.120433E-6   -1.120433E-6   -2.886193E-5   2.888367E-5   1.777769E+2   2.677769E+2   
4.162637E+3   9.004760E+1   9.004760E+1   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.849000E+3   -1.849000E+3   -2.350290E-2   2.556704E-2   -3.118213E-5   6.684714E-7   -6.684714E-7   -3.118213E-5   3.118930E-5   1.787719E+2   2.687719E+2   
4.184472E+3   9.005059E+1   9.005059E+1   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.798000E+3   -1.798000E+3   -2.441224E-2   2.609718E-2   -3.208961E-5   9.944509E-7   -9.944509E-7   -3.208961E-5   3.210501E-5   1.782250E+2   2.682250E+2   
4.206473E+3   8.996780E+1   8.996780E+1   -1.750000E+3   -1.750000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   -2.453497E-2   2.953204E-2   -3.440257E-5   -1.160386E-6   1.160386E-6   -3.440257E-5   3.442214E-5   -1.780682E+2   -8.806817E+1   
4.228446E+3   9.003301E+1   9.003301E+1   -1.700000E+3   -1.700000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   -2.575172E-2   3.000081E-2   -3.546013E-5   -5.669137E-7   5.669137E-7   -3.546013E-5   3.546466E-5   -1.790841E+2   -8.908407E+1   
4.250345E+3   9.001061E+1   9.001061E+1   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   -2.763727E-2   3.251406E-2   -3.826272E-5   -8.153915E-7   8.153915E-7   -3.826272E-5   3.827141E-5   -1.787792E+2   -8.877919E+1   
4.272179E+3   9.002200E+1   9.002200E+1   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.599000E+3   -1.599000E+3   -2.770232E-2   3.533961E-2   -4.014318E-5   -2.614546E-6   2.614546E-6   -4.014318E-5   4.022824E-5   -1.762736E+2   -8.627356E+1   
4.294313E+3   9.004681E+1   9.004681E+1   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   -2.842389E-2   3.651585E-2   -4.135536E-5   -2.849834E-6   2.849834E-6   -4.135536E-5   4.145344E-5   -1.760579E+2   -8.605793E+1   
4.316406E+3   9.001531E+1   9.001531E+1   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   -3.170044E-2   3.729081E-2   -4.388580E-5   -9.330488E-7   9.330488E-7   -4.388580E-5   4.389572E-5   -1.787820E+2   -8.878203E+1   
4.338423E+3   9.003289E+1   9.003289E+1   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   -3.347737E-2   3.980223E-2   -4.662005E-5   -1.260664E-6   1.260664E-6   -4.662005E-5   4.663709E-5   -1.784510E+2   -8.845103E+1   
4.360521E+3   9.003869E+1   9.003869E+1   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   -3.374860E-2   4.158654E-2   -4.794983E-5   -2.226592E-6   2.226592E-6   -4.794983E-5   4.800150E-5   -1.773413E+2   -8.734133E+1   
4.382343E+3   9.004199E+1   9.004199E+1   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   -3.499968E-2   4.319595E-2   -4.977151E-5   -2.353445E-6   2.353445E-6   -4.977151E-5   4.982712E-5   -1.772928E+2   -8.729279E+1   
4.404411E+3   9.001489E+1   9.001489E+1   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   -3.549608E-2   4.469375E-2   -5.105390E-5   -2.965508E-6   2.965508E-6   -5.105390E-5   5.113996E-5   -1.766757E+2   -8.667566E+1   
4.426469E+3   9.004281E+1   9.004281E+1   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   -3.723744E-2   4.730156E-2   -5.382893E-5   -3.382454E-6   3.382454E-6   -5.382893E-5   5.393510E-5   -1.764044E+2   -8.640443E+1   
4.448292E+3   9.004089E+1   9.004089E+1   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   -3.894075E-2   4.857417E-2   -5.571084E-5   -2.954629E-6   2.954629E-6   -5.571084E-5   5.578913E-5   -1.769642E+2   -8.696416E+1   
4.470347E+3   8.997561E+1   8.997561E+1   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.150000E+3   -1.150000E+3   -4.074837E-2   5.016522E-2   -5.786463E-5   -2.657841E-6   2.657841E-6   -5.786463E-5   5.792564E-5   -1.773701E+2   -8.737014E+1   
4.492376E+3   9.002551E+1   9.002551E+1   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   -4.189210E-2   5.275087E-2   -6.025574E-5   -3.502333E-6   3.502333E-6   -6.025574E-5   6.035744E-5   -1.766735E+2   -8.667346E+1   
4.514495E+3   9.001010E+1   9.001010E+1   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   -4.246581E-2   5.319327E-2   -6.089856E-5   -3.367227E-6   3.367227E-6   -6.089856E-5   6.099158E-5   -1.768352E+2   -8.683520E+1   
4.536551E+3   9.000131E+1   9.000131E+1   -1.000000E+3   -1.000000E+3   9.000000E+1   -1.000000E+3   -1.000000E+3   -4.389547E-2   5.635324E-2   -6.384050E-5   -4.375707E-6   4.375707E-6   -6.384050E-5   6.399028E-5   -1.760790E+2   -8.607901E+1   
4.558506E+3   9.002929E+1   9.002929E+1   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   -4.567367E-2   5.823879E-2   -6.616791E-5   -4.293210E-6   4.293210E-6   -6.616791E-5   6.630704E-5   -1.762876E+2   -8.628765E+1   
4.580216E+3   9.000219E+1   9.000219E+1   -9.000000E+2   -9.000000E+2   9.000000E+1   -9.000000E+2   -9.000000E+2   -4.560924E-2   5.946474E-2   -6.692652E-5   -5.142352E-6   5.142352E-6   -6.692652E-5   6.712379E-5   -1.756063E+2   -8.560627E+1   
4.602100E+3   9.002050E+1   9.002050E+1   -8.510000E+2   -8.510000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   -4.672600E-2   6.252653E-2   -6.961107E-5   -6.318078E-6   6.318078E-6   -6.961107E-5   6.989720E-5   -1.748139E+2   -8.481390E+1   
4.623774E+3   9.003881E+1   9.003881E+1   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   -4.865328E-2   6.292044E-2   -7.105915E-5   -5.150128E-6   5.150128E-6   -7.105915E-5   7.124554E-5   -1.758546E+2   -8.585464E+1   
4.645469E+3   8.998708E+1   8.998708E+1   -7.500000E+2   -7.500000E+2   9.000000E+1   -7.490000E+2   -7.490000E+2   -4.934728E-2   6.499374E-2   -7.283854E-5   -5.992290E-6   5.992290E-6   -7.283854E-5   7.308461E-5   -1.752970E+2   -8.529697E+1   
4.667347E+3   8.996621E+1   8.996621E+1   -7.010000E+2   -7.010000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   -5.226860E-2   6.619700E-2   -7.542830E-5   -4.618253E-6   4.618253E-6   -7.542830E-5   7.556955E-5   -1.764963E+2   -8.649632E+1   
4.689220E+3   9.003509E+1   9.003509E+1   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.500000E+2   -6.500000E+2   -5.232258E-2   6.852493E-2   -7.697782E-5   -6.100255E-6   6.100255E-6   -7.697782E-5   7.721916E-5   -1.754690E+2   -8.546896E+1   
4.710847E+3   9.002191E+1   9.002191E+1   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   -5.286501E-2   6.945881E-2   -7.792141E-5   -6.309600E-6   6.309600E-6   -7.792141E-5   7.817645E-5   -1.753706E+2   -8.537064E+1   
4.732786E+3   8.993020E+1   8.993020E+1   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   -5.574334E-2   7.070684E-2   -8.051375E-5   -4.996630E-6   4.996630E-6   -8.051375E-5   8.066865E-5   -1.764488E+2   -8.644882E+1   
4.754411E+3   8.997759E+1   8.997759E+1   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   -5.450633E-2   7.376189E-2   -8.173870E-5   -7.908864E-6   7.908864E-6   -8.173870E-5   8.212043E-5   -1.744734E+2   -8.447339E+1   
4.776046E+3   9.005850E+1   9.005850E+1   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   -5.771050E-2   7.476631E-2   -8.437383E-5   -6.195623E-6   6.195623E-6   -8.437383E-5   8.460100E-5   -1.758003E+2   -8.580027E+1   
4.797765E+3   8.997369E+1   8.997369E+1   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   -5.879594E-2   7.675189E-2   -8.633809E-5   -6.690916E-6   6.690916E-6   -8.633809E-5   8.659696E-5   -1.755686E+2   -8.556862E+1   
4.819406E+3   9.004339E+1   9.004339E+1   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   -6.038451E-2   7.770172E-2   -8.793883E-5   -6.136932E-6   6.136932E-6   -8.793883E-5   8.815271E-5   -1.760080E+2   -8.600801E+1   
4.841030E+3   9.001711E+1   9.001711E+1   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   -6.070540E-2   7.960198E-2   -8.937485E-5   -7.141929E-6   7.141929E-6   -8.937485E-5   8.965975E-5   -1.754312E+2   -8.543121E+1   
4.862773E+3   8.996179E+1   8.996179E+1   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   -6.301677E-2   8.099727E-2   -9.171258E-5   -6.344564E-6   6.344564E-6   -9.171258E-5   9.193177E-5   -1.760427E+2   -8.604265E+1   
4.884454E+3   9.001550E+1   9.001550E+1   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   -6.378314E-2   8.397745E-2   -9.412734E-5   -7.726098E-6   7.726098E-6   -9.412734E-5   9.444390E-5   -1.753076E+2   -8.530760E+1   
4.906145E+3   9.001931E+1   9.001931E+1   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.500000E+2   -1.500000E+2   -6.429916E-2   8.556113E-2   -9.547781E-5   -8.379792E-6   8.379792E-6   -9.547781E-5   9.584484E-5   -1.749842E+2   -8.498418E+1   
4.927816E+3   9.002130E+1   9.002130E+1   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   -6.600554E-2   8.649131E-2   -9.713859E-5   -7.725831E-6   7.725831E-6   -9.713859E-5   9.744534E-5   -1.754526E+2   -8.545260E+1   
4.949333E+3   9.004489E+1   9.004489E+1   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   -6.648475E-2   8.960896E-2   -9.946535E-5   -9.409620E-6   9.409620E-6   -9.946535E-5   9.990944E-5   -1.745958E+2   -8.459579E+1   
4.982388E+3   9.001861E+1   9.001861E+1   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.600000E+1   -4.600000E+1   -6.579509E-2   8.828297E-2   -9.817537E-5   -9.052824E-6   9.052824E-6   -9.817537E-5   9.859187E-5   -1.747316E+2   -8.473161E+1   
5.004668E+3   8.997360E+1   8.997360E+1   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   -6.657127E-2   8.778109E-2   -9.832837E-5   -8.150614E-6   8.150614E-6   -9.832837E-5   9.866560E-5   -1.752615E+2   -8.526148E+1   
5.026927E+3   8.998571E+1   8.998571E+1   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   -6.779046E-2   8.841308E-2   -9.949373E-5   -7.662045E-6   7.662045E-6   -9.949373E-5   9.978833E-5   -1.755963E+2   -8.559633E+1   
5.049185E+3   9.003188E+1   9.003188E+1   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   -6.712596E-2   8.766389E-2   -9.859497E-5   -7.663731E-6   7.663731E-6   -9.859497E-5   9.889237E-5   -1.755554E+2   -8.555537E+1   
5.071414E+3   9.001901E+1   9.001901E+1   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   -6.702717E-2   8.892051E-2   -9.935232E-5   -8.558343E-6   8.558343E-6   -9.935232E-5   9.972025E-5   -1.750766E+2   -8.507662E+1   
5.093691E+3   9.000991E+1   9.000991E+1   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   -6.704744E-2   8.851861E-2   -9.910309E-5   -8.280602E-6   8.280602E-6   -9.910309E-5   9.944844E-5   -1.752237E+2   -8.522372E+1   
5.115944E+3   9.003509E+1   9.003509E+1   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   -6.678909E-2   8.911317E-2   -9.933060E-5   -8.860388E-6   8.860388E-6   -9.933060E-5   9.972500E-5   -1.749027E+2   -8.490265E+1   
5.138225E+3   9.002331E+1   9.002331E+1   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   -6.690384E-2   8.918679E-2   -9.944950E-5   -8.823646E-6   8.823646E-6   -9.944950E-5   9.984017E-5   -1.749297E+2   -8.492972E+1   
5.160500E+3   9.001129E+1   9.001129E+1   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   -6.689033E-2   8.920337E-2   -9.945194E-5   -8.844477E-6   8.844477E-6   -9.945194E-5   9.984445E-5   -1.749179E+2   -8.491793E+1   
5.182748E+3   9.004009E+1   9.004009E+1   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   -6.661116E-2   8.896835E-2   -9.912628E-5   -8.897309E-6   8.897309E-6   -9.912628E-5   9.952477E-5   -1.748710E+2   -8.487103E+1   
5.204929E+3   8.997299E+1   8.997299E+1   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   -6.739963E-2   8.953349E-2   -9.998182E-5   -8.683607E-6   8.683607E-6   -9.998182E-5   1.003582E-4   -1.750362E+2   -8.503621E+1   
5.227181E+3   9.006121E+1   9.006121E+1   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   -6.716216E-2   8.814431E-2   -9.893024E-5   -7.951040E-6   7.951040E-6   -9.893024E-5   9.924924E-5   -1.754050E+2   -8.540501E+1   
5.249471E+3   9.001571E+1   9.001571E+1   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   -6.744993E-2   8.853947E-2   -9.936552E-5   -7.996538E-6   7.996538E-6   -9.936552E-5   9.968676E-5   -1.753990E+2   -8.539898E+1   
5.271746E+3   8.999041E+1   8.999041E+1   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   -6.578772E-2   8.886036E-2   -9.854686E-5   -9.435756E-6   9.435756E-6   -9.854686E-5   9.899756E-5   -1.745307E+2   -8.453066E+1   
5.293993E+3   8.999490E+1   8.999490E+1   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   -6.625466E-2   8.929725E-2   -9.912008E-5   -9.376015E-6   9.376015E-6   -9.912008E-5   9.956254E-5   -1.745963E+2   -8.459633E+1   
5.316235E+3   9.002700E+1   9.002700E+1   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   -6.743950E-2   8.955436E-2   -1.000201E-4   -8.667761E-6   8.667761E-6   -1.000201E-4   1.003949E-4   -1.750471E+2   -8.504711E+1   
5.338418E+3   9.001391E+1   9.001391E+1   -1.500000E+1   -1.500000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   -6.663018E-2   8.948624E-2   -9.947533E-5   -9.221826E-6   9.221826E-6   -9.947533E-5   9.990187E-5   -1.747036E+2   -8.470355E+1   
5.359697E+3   9.001339E+1   9.001339E+1   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   -6.793282E-2   8.971145E-2   -1.004274E-4   -8.405593E-6   8.405593E-6   -1.004274E-4   1.007785E-4   -1.752156E+2   -8.521560E+1   
5.381876E+3   8.999490E+1   8.999490E+1   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   -6.701735E-2   9.061034E-2   -1.004468E-4   -9.670368E-6   9.670368E-6   -1.004468E-4   1.009112E-4   -1.745009E+2   -8.450088E+1   
5.404075E+3   9.003671E+1   9.003671E+1   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   -6.736955E-2   9.043548E-2   -1.005507E-4   -9.295550E-6   9.295550E-6   -1.005507E-4   1.009794E-4   -1.747182E+2   -8.471822E+1   
5.426155E+3   9.000881E+1   9.000881E+1   -7.000000E+0   -7.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   -6.686581E-2   8.948623E-2   -9.962100E-5   -9.047542E-6   9.047542E-6   -9.962100E-5   1.000310E-4   -1.748107E+2   -8.481065E+1   
5.447236E+3   9.001611E+1   9.001611E+1   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   -6.743030E-2   9.123192E-2   -1.011069E-4   -9.771310E-6   9.771310E-6   -1.011069E-4   1.015780E-4   -1.744799E+2   -8.447989E+1   
5.469312E+3   8.999401E+1   8.999401E+1   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   -6.698484E-2   9.038392E-2   -1.002793E-4   -9.546391E-6   9.546391E-6   -1.002793E-4   1.007326E-4   -1.745619E+2   -8.456194E+1   
5.491401E+3   9.003939E+1   9.003939E+1   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   -6.566869E-2   9.032073E-2   -9.942439E-5   -1.047853E-5   1.047853E-5   -9.942439E-5   9.997504E-5   -1.739837E+2   -8.398369E+1   
5.513419E+3   9.000631E+1   9.000631E+1   0.000000E+0   0.000000E+0   9.000000E+1   0.000000E+0   0.000000E+0   -6.757019E-2   8.957340E-2   -1.001133E-4   -8.583543E-6   8.583543E-6   -1.001133E-4   1.004806E-4   -1.750995E+2   -8.509954E+1   
5.535602E+3   9.005499E+1   9.005499E+1   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   -6.876731E-2   9.000472E-2   -1.011343E-4   -7.980110E-6   7.980110E-6   -1.011343E-4   1.014486E-4   -1.754884E+2   -8.548836E+1   
5.557103E+3   8.999890E+1   8.999890E+1   3.000000E+0   3.000000E+0   9.000000E+1   3.000000E+0   3.000000E+0   -6.829484E-2   9.122638E-2   -1.016378E-4   -9.128246E-6   9.128246E-6   -1.016378E-4   1.020469E-4   -1.748679E+2   -8.486795E+1   
5.578763E+3   9.004171E+1   9.004171E+1   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   -6.798621E-2   9.068401E-2   -1.010938E-4   -9.001934E-6   9.001934E-6   -1.010938E-4   1.014938E-4   -1.749115E+2   -8.491150E+1   
5.600302E+3   9.002609E+1   9.002609E+1   7.000000E+0   7.000000E+0   9.000000E+1   8.000000E+0   8.000000E+0   -6.782054E-2   8.965680E-2   -1.003224E-4   -8.452905E-6   8.452905E-6   -1.003224E-4   1.006778E-4   -1.751838E+2   -8.518378E+1   
5.621975E+3   9.005441E+1   9.005441E+1   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   -7.035770E-2   9.012805E-2   -1.021979E-4   -6.884432E-6   6.884432E-6   -1.021979E-4   1.024295E-4   -1.761462E+2   -8.614616E+1   
5.643832E+3   9.004699E+1   9.004699E+1   1.000000E+1   1.000000E+1   9.000000E+1   1.100000E+1   1.100000E+1   -6.926982E-2   9.003295E-2   -1.014634E-4   -7.626891E-6   7.626891E-6   -1.014634E-4   1.017496E-4   -1.757012E+2   -8.570122E+1   
5.665662E+3   9.005929E+1   9.005929E+1   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   -6.790399E-2   9.077906E-2   -1.011049E-4   -9.124884E-6   9.124884E-6   -1.011049E-4   1.015158E-4   -1.748429E+2   -8.484293E+1   
5.687504E+3   9.006539E+1   9.006539E+1   1.500000E+1   1.500000E+1   9.000000E+1   1.500000E+1   1.500000E+1   -6.792912E-2   9.193512E-2   -1.018733E-4   -9.862097E-6   9.862097E-6   -1.018733E-4   1.023496E-4   -1.744706E+2   -8.447057E+1   
5.709566E+3   9.001360E+1   9.001360E+1   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   -6.767388E-2   9.031336E-2   -1.006593E-4   -8.990618E-6   8.990618E-6   -1.006593E-4   1.010600E-4   -1.748960E+2   -8.489604E+1   
5.731434E+3   9.001339E+1   9.001339E+1   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   -6.821202E-2   9.087722E-2   -1.013592E-4   -8.961236E-6   8.961236E-6   -1.013592E-4   1.017546E-4   -1.749476E+2   -8.494758E+1   
5.753302E+3   8.996249E+1   8.996249E+1   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   -6.854949E-2   9.059807E-2   -1.013861E-4   -8.529132E-6   8.529132E-6   -1.013861E-4   1.017442E-4   -1.751913E+2   -8.519130E+1   
5.775159E+3   9.003369E+1   9.003369E+1   2.200000E+1   2.200000E+1   9.000000E+1   2.300000E+1   2.300000E+1   -6.825863E-2   9.120490E-2   -1.016015E-4   -9.140990E-6   9.140990E-6   -1.016015E-4   1.020118E-4   -1.748590E+2   -8.485899E+1   
5.797021E+3   9.003289E+1   9.003289E+1   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   -6.893848E-2   9.124910E-2   -1.020506E-4   -8.667048E-6   8.667048E-6   -1.020506E-4   1.024179E-4   -1.751456E+2   -8.514558E+1   
5.818862E+3   9.003591E+1   9.003591E+1   2.600000E+1   2.600000E+1   9.000000E+1   2.700000E+1   2.700000E+1   -6.899187E-2   9.177618E-2   -1.024269E-4   -8.972147E-6   8.972147E-6   -1.024269E-4   1.028191E-4   -1.749939E+2   -8.499392E+1   
5.840769E+3   9.001129E+1   9.001129E+1   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   -6.902377E-2   9.104722E-2   -1.019718E-4   -8.471978E-6   8.471978E-6   -1.019718E-4   1.023231E-4   -1.752507E+2   -8.525068E+1   
5.862635E+3   9.000961E+1   9.000961E+1   3.000000E+1   3.000000E+1   9.000000E+1   3.100000E+1   3.100000E+1   -6.923178E-2   9.048334E-2   -1.017332E-4   -7.949478E-6   7.949478E-6   -1.017332E-4   1.020433E-4   -1.755320E+2   -8.553196E+1   
5.884570E+3   9.006179E+1   9.006179E+1   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   -6.922443E-2   9.087236E-2   -1.019820E-4   -8.209242E-6   8.209242E-6   -1.019820E-4   1.023119E-4   -1.753978E+2   -8.539779E+1   
5.906445E+3   9.004839E+1   9.004839E+1   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   -6.919434E-2   9.147303E-2   -1.023546E-4   -8.624198E-6   8.624198E-6   -1.023546E-4   1.027173E-4   -1.751837E+2   -8.518375E+1   
5.928319E+3   9.000891E+1   9.000891E+1   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   -6.803346E-2   9.261254E-2   -1.023790E-4   -1.022780E-5   1.022780E-5   -1.023790E-4   1.028886E-4   -1.742950E+2   -8.429500E+1   
5.950188E+3   9.003469E+1   9.003469E+1   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   -6.879859E-2   9.183875E-2   -1.023481E-4   -9.156008E-6   9.156008E-6   -1.023481E-4   1.027568E-4   -1.748880E+2   -8.488796E+1   
5.972023E+3   8.997521E+1   8.997521E+1   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   -6.844822E-2   9.307027E-2   -1.029336E-4   -1.022028E-5   1.022028E-5   -1.029336E-4   1.034397E-4   -1.743297E+2   -8.432968E+1   
5.993898E+3   8.997720E+1   8.997720E+1   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   -6.858813E-2   9.142765E-2   -1.019503E-4   -9.042902E-6   9.042902E-6   -1.019503E-4   1.023505E-4   -1.749312E+2   -8.493118E+1   
6.015829E+3   9.000131E+1   9.000131E+1   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   -6.862065E-2   9.194062E-2   -1.023044E-4   -9.354219E-6   9.354219E-6   -1.023044E-4   1.027312E-4   -1.747757E+2   -8.477568E+1   
6.037662E+3   8.995172E+1   8.995172E+1   4.600000E+1   4.600000E+1   9.000000E+1   4.700000E+1   4.700000E+1   -6.892252E-2   9.204310E-2   -1.025578E-4   -9.197942E-6   9.197942E-6   -1.025578E-4   1.029695E-4   -1.748751E+2   -8.487512E+1   
6.059575E+3   8.999410E+1   8.999410E+1   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   -6.922994E-2   9.112698E-2   -1.021512E-4   -8.371635E-6   8.371635E-6   -1.021512E-4   1.024937E-4   -1.753149E+2   -8.531489E+1   
6.093454E+3   9.007650E+1   9.007650E+1   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   -6.894892E-2   9.382013E-2   -1.037315E-4   -1.034019E-5   1.034019E-5   -1.037315E-4   1.042456E-4   -1.743074E+2   -8.430743E+1   
6.115976E+3   9.002331E+1   9.002331E+1   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   -7.100197E-2   9.619118E-2   -1.065450E-4   -1.037181E-5   1.037181E-5   -1.065450E-4   1.070487E-4   -1.744400E+2   -8.443996E+1   
6.138088E+3   9.005050E+1   9.005050E+1   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   -7.204324E-2   9.692322E-2   -1.076656E-4   -1.008024E-5   1.008024E-5   -1.076656E-4   1.081364E-4   -1.746512E+2   -8.465125E+1   
6.160257E+3   9.007299E+1   9.007299E+1   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   -7.405763E-2   9.826086E-2   -1.097821E-4   -9.464855E-6   9.464855E-6   -1.097821E-4   1.101894E-4   -1.750724E+2   -8.507244E+1   
6.183075E+3   8.998531E+1   8.998531E+1   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   -7.499763E-2   1.008269E-1   -1.120345E-4   -1.044719E-5   1.044719E-5   -1.120345E-4   1.125206E-4   -1.746726E+2   -8.467259E+1   
6.205450E+3   8.994641E+1   8.994641E+1   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   -7.610639E-2   1.009128E-1   -1.127759E-4   -9.683263E-6   9.683263E-6   -1.127759E-4   1.131909E-4   -1.750925E+2   -8.509246E+1   
6.227739E+3   9.004958E+1   9.004958E+1   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   -7.667396E-2   1.025271E-1   -1.141783E-4   -1.031890E-5   1.031890E-5   -1.141783E-4   1.146436E-4   -1.748359E+2   -8.483590E+1   
6.250620E+3   9.000790E+1   9.000790E+1   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   -7.874174E-2   1.052342E-1   -1.172198E-4   -1.055933E-5   1.055933E-5   -1.172198E-4   1.176944E-4   -1.748526E+2   -8.485260E+1   
6.272755E+3   9.004891E+1   9.004891E+1   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   -8.003948E-2   1.058828E-1   -1.184445E-4   -1.002349E-5   1.002349E-5   -1.184445E-4   1.188679E-4   -1.751628E+2   -8.516281E+1   
6.295331E+3   9.006021E+1   9.006021E+1   5.480000E+2   5.480000E+2   9.000000E+1   5.480000E+2   5.480000E+2   -8.048187E-2   1.073161E-1   -1.196515E-4   -1.063337E-5   1.063337E-5   -1.196515E-4   1.201231E-4   -1.749215E+2   -8.492149E+1   
6.318620E+3   9.002929E+1   9.002929E+1   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   -8.141206E-2   1.094097E-1   -1.215901E-4   -1.131408E-5   1.131408E-5   -1.215901E-4   1.221154E-4   -1.746839E+2   -8.468388E+1   
6.341226E+3   9.003781E+1   9.003781E+1   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   -8.185138E-2   1.113357E-1   -1.231161E-4   -1.224833E-5   1.224833E-5   -1.231161E-4   1.237239E-4   -1.743186E+2   -8.431857E+1   
6.364104E+3   9.007711E+1   9.007711E+1   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   -8.265702E-2   1.126733E-1   -1.244854E-4   -1.252695E-5   1.252695E-5   -1.244854E-4   1.251141E-4   -1.742537E+2   -8.425368E+1   
6.387565E+3   9.003771E+1   9.003771E+1   7.480000E+2   7.480000E+2   9.000000E+1   7.480000E+2   7.480000E+2   -8.445114E-2   1.143251E-1   -1.266704E-4   -1.227985E-5   1.227985E-5   -1.266704E-4   1.272642E-4   -1.744629E+2   -8.446286E+1   
6.410192E+3   9.004269E+1   9.004269E+1   7.980000E+2   7.980000E+2   9.000000E+1   7.980000E+2   7.980000E+2   -8.513407E-2   1.171059E-1   -1.289037E-4   -1.359272E-5   1.359272E-5   -1.289037E-4   1.296184E-4   -1.739805E+2   -8.398048E+1   
6.432727E+3   9.000210E+1   9.000210E+1   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   -8.528009E-2   1.179643E-1   -1.295530E-4   -1.404593E-5   1.404593E-5   -1.295530E-4   1.303122E-4   -1.738123E+2   -8.381225E+1   
6.455974E+3   9.002029E+1   9.002029E+1   8.980000E+2   8.980000E+2   9.000000E+1   8.980000E+2   8.980000E+2   -8.766265E-2   1.185245E-1   -1.313909E-4   -1.264995E-5   1.264995E-5   -1.313909E-4   1.319984E-4   -1.745007E+2   -8.450067E+1   
6.478551E+3   9.001171E+1   9.001171E+1   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   -8.841981E-2   1.207224E-1   -1.332905E-4   -1.352683E-5   1.352683E-5   -1.332905E-4   1.339751E-4   -1.742052E+2   -8.420524E+1   
6.501119E+3   9.003301E+1   9.003301E+1   9.980000E+2   9.980000E+2   9.000000E+1   9.980000E+2   9.980000E+2   -8.981942E-2   1.221140E-1   -1.350621E-4   -1.340143E-5   1.340143E-5   -1.350621E-4   1.357253E-4   -1.743334E+2   -8.433342E+1   
6.524662E+3   9.007491E+1   9.007491E+1   1.048000E+3   1.048000E+3   9.000000E+1   1.048000E+3   1.048000E+3   -9.056065E-2   1.233184E-1   -1.363048E-4   -1.364064E-5   1.364064E-5   -1.363048E-4   1.369857E-4   -1.742852E+2   -8.428518E+1   
6.547448E+3   9.003521E+1   9.003521E+1   1.098000E+3   1.098000E+3   9.000000E+1   1.098000E+3   1.098000E+3   -9.174976E-2   1.253089E-1   -1.383364E-4   -1.406245E-5   1.406245E-5   -1.383364E-4   1.390493E-4   -1.741956E+2   -8.419559E+1   
6.570284E+3   9.006078E+1   9.006078E+1   1.148000E+3   1.148000E+3   9.000000E+1   1.148000E+3   1.148000E+3   -9.271442E-2   1.272448E-1   -1.401936E-4   -1.461457E-5   1.461457E-5   -1.401936E-4   1.409533E-4   -1.740487E+2   -8.404866E+1   
6.593584E+3   8.998651E+1   8.998651E+1   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   -9.453375E-2   1.281406E-1   -1.419018E-4   -1.385461E-5   1.385461E-5   -1.419018E-4   1.425766E-4   -1.744236E+2   -8.442359E+1   
6.616471E+3   9.003839E+1   9.003839E+1   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   -9.417361E-2   1.309159E-1   -1.434866E-4   -1.593537E-5   1.593537E-5   -1.434866E-4   1.443688E-4   -1.736628E+2   -8.366280E+1   
6.639463E+3   9.006329E+1   9.006329E+1   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   -9.596530E-2   1.320528E-1   -1.453348E-4   -1.535349E-5   1.535349E-5   -1.453348E-4   1.461436E-4   -1.739695E+2   -8.396952E+1   
6.663064E+3   9.006100E+1   9.006100E+1   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   -9.738582E-2   1.339464E-1   -1.474463E-4   -1.554077E-5   1.554077E-5   -1.474463E-4   1.482630E-4   -1.739833E+2   -8.398327E+1   
6.685646E+3   9.004559E+1   9.004559E+1   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   -9.799272E-2   1.345004E-1   -1.481824E-4   -1.545411E-5   1.545411E-5   -1.481824E-4   1.489861E-4   -1.740461E+2   -8.404608E+1   
6.708427E+3   9.002661E+1   9.002661E+1   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   -9.886277E-2   1.359896E-1   -1.496902E-4   -1.578418E-5   1.578418E-5   -1.496902E-4   1.505200E-4   -1.739807E+2   -8.398065E+1   
6.731470E+3   9.000839E+1   9.000839E+1   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   -9.949476E-2   1.373462E-1   -1.509645E-4   -1.620366E-5   1.620366E-5   -1.509645E-4   1.518316E-4   -1.738737E+2   -8.387365E+1   
6.754042E+3   9.003680E+1   9.003680E+1   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   -1.009484E-1   1.384145E-1   -1.525589E-4   -1.582693E-5   1.582693E-5   -1.525589E-4   1.533776E-4   -1.740771E+2   -8.407715E+1   
6.776578E+3   9.000741E+1   9.000741E+1   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   -1.030161E-1   1.405792E-1   -1.552471E-4   -1.571277E-5   1.571277E-5   -1.552471E-4   1.560403E-4   -1.742207E+2   -8.422070E+1   
6.799610E+3   9.003201E+1   9.003201E+1   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   -1.032554E-1   1.422469E-1   -1.564813E-4   -1.662609E-5   1.662609E-5   -1.564813E-4   1.573620E-4   -1.739351E+2   -8.393509E+1   
6.822190E+3   9.004269E+1   9.004269E+1   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   -1.038758E-1   1.438024E-1   -1.578778E-4   -1.718418E-5   1.718418E-5   -1.578778E-4   1.588103E-4   -1.737881E+2   -8.378810E+1   
6.844770E+3   9.003860E+1   9.003860E+1   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   -1.046630E-1   1.439146E-1   -1.584376E-4   -1.667532E-5   1.667532E-5   -1.584376E-4   1.593128E-4   -1.739918E+2   -8.399182E+1   
6.867549E+3   9.002691E+1   9.002691E+1   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   -1.062068E-1   1.467580E-1   -1.612439E-4   -1.739240E-5   1.739240E-5   -1.612439E-4   1.621792E-4   -1.738437E+2   -8.384365E+1   
6.890127E+3   9.002340E+1   9.002340E+1   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   -1.084531E-1   1.487325E-1   -1.639187E-4   -1.702184E-5   1.702184E-5   -1.639187E-4   1.648001E-4   -1.740715E+2   -8.407147E+1   
6.912611E+3   8.999420E+1   8.999420E+1   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   -1.113087E-1   1.505076E-1   -1.668403E-4   -1.607024E-5   1.607024E-5   -1.668403E-4   1.676125E-4   -1.744982E+2   -8.449818E+1   
6.935698E+3   8.995400E+1   8.995400E+1   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   -1.093428E-1   1.519538E-1   -1.665668E-4   -1.846976E-5   1.846976E-5   -1.665668E-4   1.675877E-4   -1.736726E+2   -8.367260E+1   
6.958219E+3   9.002041E+1   9.002041E+1   1.998000E+3   1.998000E+3   9.000000E+1   1.999000E+3   1.999000E+3   -1.108989E-1   1.543198E-1   -1.690697E-4   -1.886569E-5   1.886569E-5   -1.690697E-4   1.701190E-4   -1.736330E+2   -8.363297E+1   
6.996117E+3   9.004351E+1   9.004351E+1   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   -1.219446E-1   1.702332E-1   -1.862629E-4   -2.109960E-5   2.109960E-5   -1.862629E-4   1.874542E-4   -1.735372E+2   -8.353716E+1   
7.023020E+3   9.001840E+1   9.001840E+1   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   -1.358215E-1   1.890774E-1   -2.071153E-4   -2.315569E-5   2.315569E-5   -2.071153E-4   2.084057E-4   -1.736208E+2   -8.362077E+1   
7.048969E+3   8.999539E+1   8.999539E+1   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -1.483000E-1   2.084068E-1   -2.274191E-4   -2.656325E-5   2.656325E-5   -2.274191E-4   2.289652E-4   -1.733379E+2   -8.333787E+1   
7.074904E+3   9.000021E+1   9.000021E+1   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -1.602735E-1   2.246043E-1   -2.453709E-4   -2.829670E-5   2.829670E-5   -2.453709E-4   2.469971E-4   -1.734216E+2   -8.342159E+1   
7.101389E+3   9.006329E+1   9.006329E+1   4.498000E+3   4.498000E+3   9.000000E+1   4.499000E+3   4.499000E+3   -1.668554E-1   2.371208E-1   -2.575921E-4   -3.161145E-5   3.161145E-5   -2.575921E-4   2.595245E-4   -1.730037E+2   -8.300370E+1   
7.127483E+3   9.002731E+1   9.002731E+1   4.997000E+3   4.997000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -1.678923E-1   2.422816E-1   -2.615943E-4   -3.421851E-5   3.421851E-5   -2.615943E-4   2.638229E-4   -1.725476E+2   -8.254759E+1   
7.153214E+3   9.001379E+1   9.001379E+1   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -1.608913E-1   2.358801E-1   -2.530968E-4   -3.521154E-5   3.521154E-5   -2.530968E-4   2.555344E-4   -1.720797E+2   -8.207969E+1   
7.179579E+3   8.997759E+1   8.997759E+1   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -1.450369E-1   2.199698E-1   -2.329326E-4   -3.653628E-5   3.653628E-5   -2.329326E-4   2.357806E-4   -1.710856E+2   -8.108559E+1   
7.205482E+3   9.000839E+1   9.000839E+1   6.497000E+3   6.497000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -1.284296E-1   2.005744E-1   -2.100332E-4   -3.613937E-5   3.613937E-5   -2.100332E-4   2.131197E-4   -1.702370E+2   -8.023700E+1   
7.231627E+3   8.998019E+1   8.998019E+1   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -1.205144E-1   1.919725E-1   -1.995372E-4   -3.637001E-5   3.637001E-5   -1.995372E-4   2.028248E-4   -1.696700E+2   -7.967000E+1   
7.257521E+3   9.005239E+1   9.005239E+1   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -1.132544E-1   1.863130E-1   -1.913629E-4   -3.803971E-5   3.803971E-5   -1.913629E-4   1.951071E-4   -1.687571E+2   -7.875712E+1   
7.283356E+3   9.002569E+1   9.002569E+1   7.999000E+3   7.999000E+3   9.000000E+1   8.000000E+3   8.000000E+3   -1.164058E-1   1.926480E-1   -1.974371E-4   -3.985050E-5   3.985050E-5   -1.974371E-4   2.014187E-4   -1.685888E+2   -7.858879E+1   
7.309758E+3   9.002761E+1   9.002761E+1   8.498000E+3   8.498000E+3   9.000000E+1   8.499000E+3   8.499000E+3   -1.229251E-1   2.045124E-1   -2.091948E-4   -4.278520E-5   4.278520E-5   -2.091948E-4   2.135253E-4   -1.684411E+2   -7.844109E+1   
7.336115E+3   8.997280E+1   8.997280E+1   8.998000E+3   8.998000E+3   9.000000E+1   8.999000E+3   8.999000E+3   -1.317694E-1   2.166050E-1   -2.225385E-4   -4.414948E-5   4.414948E-5   -2.225385E-4   2.268756E-4   -1.687788E+2   -7.877878E+1   
7.362472E+3   8.997241E+1   8.997241E+1   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -1.482177E-1   2.366072E-1   -2.457349E-4   -4.506068E-5   4.506068E-5   -2.457349E-4   2.498322E-4   -1.696090E+2   -7.960905E+1   
7.387947E+3   9.001260E+1   9.001260E+1   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -1.590033E-1   2.543814E-1   -2.639792E-4   -4.870360E-5   4.870360E-5   -2.639792E-4   2.684345E-4   -1.695466E+2   -7.954660E+1   
@@END Data.
@Time at end of measurement: 15:03:08
@NO Instrument  Changes.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -9499.000      -9999.000      250.000        Coercive Field: Field at which M//H changes sign
Ms  emu                                 3.344E-4       -4.020E-4      3.682E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -1.001E-4      1.348E-4       1.174E-4       Remanent Magnetization: M at H=0        
S                                       0.299          0.335          0.317          Squareness: Mr/Ms                       
S*                                      1.221          1.296          1.259          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
