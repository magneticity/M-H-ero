@Filename: c:\vsm-lv\Will\data\AJA335e-FePtFeRh_1030nm_Tann_6\AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_140deg.VHD
@Measurement Controlfilename: C:\vsm-lv\Will\Recipes\10kOe OoP loop 140deg.VHC
@Signal Manipulation filename: c:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA335e-FePtFeRh_1030nm_Tann_6
@Date: 12 November 2019    (2019-12-11)
@Time: 10:46:33
@Test ID: AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_140deg
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 90.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Sample Temperature to 140.1478 [degC] and wait 60.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Applied Field to 9999.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 3:      Set Auto Range Signal to 11.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 5
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 5.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 10000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To: 50.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: 50.0000 [Oe] To: -50.0000 [Oe] Min Stepsize/Sweeprate =  2.0000 [Oe] Max Stepsize/Sweeprate =  2.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -50.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -10000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 4 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 10 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.706
@Y Coils Correction Factor: 0.964
@Sample Shape Correction Factor: 0.919
@Coil Angle Alpha: 42.300
@Coil Angle Beta: -47.320
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
15000.000000   1.000000
15249.000000   1.000524
15499.000000   1.000702
15750.000000   1.001233
16000.000000   1.001406
16250.000000   1.001585
16499.000000   1.001758
16749.000000   1.001937
16999.000000   1.002110
17249.000000   1.001937
17499.000000   1.002289
17749.000000   1.002289
17999.000000   1.002289
18249.000000   1.002462
18499.000000   1.002462
18748.000000   1.002462
18999.000000   1.002462
19249.000000   1.002462
19499.000000   1.002642
19749.000000   1.002642
19999.000000   1.002462
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = No
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 25 October 2019  12:02:56
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 5
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 10:46:33
@@Data
New Section: Section 0: 
3.211500E+1   1.400683E+2   1.400683E+2   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -8.289389E-2   1.968182E-1   -1.794345E-4   -6.736329E-5   6.736329E-5   -1.794345E-4   1.916626E-4   -1.594229E+2   -6.942286E+1   
5.745900E+1   1.399645E+2   1.399645E+2   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -7.210197E-2   1.793455E-1   -1.613827E-4   -6.392219E-5   6.392219E-5   -1.613827E-4   1.735811E-4   -1.583919E+2   -6.839194E+1   
8.296200E+1   1.400356E+2   1.400356E+2   8.998000E+3   8.998000E+3   9.000000E+1   8.998000E+3   8.998000E+3   -6.192996E-2   1.633185E-1   -1.446556E-4   -6.096772E-5   6.096772E-5   -1.446556E-4   1.569787E-4   -1.571461E+2   -6.714613E+1   
1.081490E+2   1.400355E+2   1.400355E+2   8.498000E+3   8.498000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -5.165281E-2   1.458088E-1   -1.268979E-4   -5.712165E-5   5.712165E-5   -1.268979E-4   1.391616E-4   -1.557657E+2   -6.576565E+1   
1.341160E+2   1.400190E+2   1.400190E+2   7.999000E+3   7.999000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -4.123972E-2   1.280270E-1   -1.088789E-4   -5.319823E-5   5.319823E-5   -1.088789E-4   1.211803E-4   -1.539599E+2   -6.395987E+1   
1.599080E+2   1.400873E+2   1.400873E+2   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -3.330604E-2   1.121955E-1   -9.366310E-5   -4.871609E-5   4.871609E-5   -9.366310E-5   1.055748E-4   -1.525201E+2   -6.252014E+1   
1.848070E+2   1.399914E+2   1.399914E+2   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -1.728311E-2   9.167973E-2   -7.039526E-5   -4.715450E-5   4.715450E-5   -7.039526E-5   8.472921E-5   -1.461837E+2   -5.618372E+1   
2.101900E+2   1.400868E+2   1.400868E+2   6.497000E+3   6.497000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -9.935073E-3   7.673424E-2   -5.611852E-5   -4.281839E-5   4.281839E-5   -5.611852E-5   7.058827E-5   -1.426564E+2   -5.265639E+1   
2.357430E+2   1.400149E+2   1.400149E+2   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -4.686290E-4   6.285802E-2   -4.122849E-5   -4.074819E-5   4.074819E-5   -4.122849E-5   5.796726E-5   -1.353357E+2   -4.533569E+1   
2.611030E+2   1.400006E+2   1.400006E+2   5.498000E+3   5.498000E+3   9.000000E+1   5.498000E+3   5.498000E+3   6.048909E-3   4.668503E-2   -2.666575E-5   -3.499532E-5   3.499532E-5   -2.666575E-5   4.399698E-5   -1.273067E+2   -3.730669E+1   
2.867390E+2   1.400931E+2   1.400931E+2   4.997000E+3   4.997000E+3   9.000000E+1   4.998000E+3   4.998000E+3   1.873929E-2   2.961409E-2   -7.701837E-6   -3.322102E-5   3.322102E-5   -7.701837E-6   3.410212E-5   -1.030526E+2   -1.305265E+1   
3.119760E+2   1.400145E+2   1.400145E+2   4.498000E+3   4.498000E+3   9.000000E+1   4.498000E+3   4.498000E+3   2.661319E-2   1.334217E-2   7.763903E-6   -2.840668E-5   2.840668E-5   7.763903E-6   2.944856E-5   -7.471367E+1   1.528633E+1   
3.382160E+2   1.400359E+2   1.400359E+2   3.999000E+3   3.999000E+3   9.000000E+1   3.999000E+3   3.999000E+3   3.515723E-2   -3.879411E-4   2.198850E-5   -2.574975E-5   2.574975E-5   2.198850E-5   3.386066E-5   -4.950497E+1   4.049503E+1   
3.636630E+2   1.400235E+2   1.400235E+2   3.498000E+3   3.498000E+3   9.000000E+1   3.498000E+3   3.498000E+3   4.717777E-2   -1.724582E-2   4.039952E-5   -2.361932E-5   2.361932E-5   4.039952E-5   4.679737E-5   -3.031241E+1   5.968759E+1   
3.885910E+2   1.400300E+2   1.400300E+2   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   5.803018E-2   -3.586346E-2   5.923446E-5   -1.947440E-5   1.947440E-5   5.923446E-5   6.235362E-5   -1.819922E+1   7.180078E+1   
4.141450E+2   1.400985E+2   1.400985E+2   2.498000E+3   2.498000E+3   9.000000E+1   2.498000E+3   2.498000E+3   6.695322E-2   -5.217916E-2   7.537735E-5   -1.540742E-5   1.540742E-5   7.537735E-5   7.693590E-5   -1.155234E+1   7.844766E+1   
4.399610E+2   1.400612E+2   1.400612E+2   1.999000E+3   1.999000E+3   9.000000E+1   1.999000E+3   1.999000E+3   7.814027E-2   -6.897224E-2   9.323086E-5   -1.270287E-5   1.270287E-5   9.323086E-5   9.409227E-5   -7.758876E+0   8.224112E+1   
4.737450E+2   1.400536E+2   1.400536E+2   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   7.977916E-2   -7.061388E-2   9.531328E-5   -1.284178E-5   1.284178E-5   9.531328E-5   9.617449E-5   -7.673387E+0   8.232661E+1   
4.960340E+2   1.400242E+2   1.400242E+2   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   8.183635E-2   -7.236781E-2   9.772745E-5   -1.321668E-5   1.321668E-5   9.772745E-5   9.861711E-5   -7.701963E+0   8.229804E+1   
5.182610E+2   1.400529E+2   1.400529E+2   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   8.307150E-2   -7.464729E-2   9.997567E-5   -1.263997E-5   1.263997E-5   9.997567E-5   1.007715E-4   -7.205702E+0   8.279430E+1   
5.404920E+2   1.400172E+2   1.400172E+2   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   8.278848E-2   -7.595928E-2   1.006552E-4   -1.157290E-5   1.157290E-5   1.006552E-4   1.013183E-4   -6.558822E+0   8.344118E+1   
5.627230E+2   1.399562E+2   1.399562E+2   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   8.508760E-2   -7.779636E-2   1.032731E-4   -1.207237E-5   1.207237E-5   1.032731E-4   1.039763E-4   -6.667475E+0   8.333252E+1   
5.849970E+2   1.400610E+2   1.400610E+2   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   8.486763E-2   -7.917109E-2   1.040324E-4   -1.101091E-5   1.101091E-5   1.040324E-4   1.046135E-4   -6.041757E+0   8.395824E+1   
6.072830E+2   1.400149E+2   1.400149E+2   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   8.718236E-2   -8.138231E-2   1.069036E-4   -1.127733E-5   1.127733E-5   1.069036E-4   1.074968E-4   -6.021895E+0   8.397810E+1   
6.296040E+2   1.399997E+2   1.399997E+2   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   8.788479E-2   -8.297010E-2   1.083720E-4   -1.075882E-5   1.075882E-5   1.083720E-4   1.089048E-4   -5.669557E+0   8.433044E+1   
6.518440E+2   1.400108E+2   1.400108E+2   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   8.890762E-2   -8.386241E-2   1.095855E-4   -1.093196E-5   1.093196E-5   1.095855E-4   1.101295E-4   -5.696826E+0   8.430317E+1   
6.740480E+2   1.400275E+2   1.400275E+2   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   9.064364E-2   -8.566573E-2   1.118333E-4   -1.103701E-5   1.103701E-5   1.118333E-4   1.123766E-4   -5.636361E+0   8.436364E+1   
6.962720E+2   1.400894E+2   1.400894E+2   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   9.150375E-2   -8.823022E-2   1.140353E-4   -9.996590E-6   9.996590E-6   1.140353E-4   1.144726E-4   -5.009869E+0   8.499013E+1   
7.185010E+2   1.400649E+2   1.400649E+2   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   9.204881E-2   -8.955003E-2   1.152319E-4   -9.536883E-6   9.536883E-6   1.152319E-4   1.156258E-4   -4.731162E+0   8.526884E+1   
7.407910E+2   1.400274E+2   1.400274E+2   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   9.450480E-2   -9.164670E-2   1.181158E-4   -9.982666E-6   9.982666E-6   1.181158E-4   1.185369E-4   -4.830925E+0   8.516908E+1   
7.630810E+2   1.400102E+2   1.400102E+2   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   9.450201E-2   -9.365601E-2   1.194227E-4   -8.666971E-6   8.666971E-6   1.194227E-4   1.197368E-4   -4.150900E+0   8.584910E+1   
7.853310E+2   1.401042E+2   1.401042E+2   1.248000E+3   1.248000E+3   9.000000E+1   1.248000E+3   1.248000E+3   9.588523E-2   -9.597532E-2   1.217884E-4   -8.173743E-6   8.173743E-6   1.217884E-4   1.220624E-4   -3.839607E+0   8.616039E+1   
8.075500E+2   1.400088E+2   1.400088E+2   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   9.730408E-2   -9.810942E-2   1.240556E-4   -7.827951E-6   7.827951E-6   1.240556E-4   1.243023E-4   -3.610598E+0   8.638940E+1   
8.298700E+2   1.400615E+2   1.400615E+2   1.147000E+3   1.147000E+3   9.000000E+1   1.148000E+3   1.148000E+3   9.834719E-2   -9.789882E-2   1.245633E-4   -8.737150E-6   8.737150E-6   1.245633E-4   1.248693E-4   -4.012284E+0   8.598772E+1   
8.521120E+2   1.400956E+2   1.400956E+2   1.097000E+3   1.097000E+3   9.000000E+1   1.098000E+3   1.098000E+3   9.908137E-2   -1.000090E-1   1.263915E-4   -7.900622E-6   7.900622E-6   1.263915E-4   1.266382E-4   -3.576855E+0   8.642315E+1   
8.744420E+2   1.400858E+2   1.400858E+2   1.047000E+3   1.047000E+3   9.000000E+1   1.048000E+3   1.048000E+3   9.930808E-2   -1.011570E-1   1.272794E-4   -7.317763E-6   7.317763E-6   1.272794E-4   1.274896E-4   -3.290524E+0   8.670948E+1   
8.965330E+2   1.400964E+2   1.400964E+2   9.980000E+2   9.980000E+2   9.000000E+1   9.990000E+2   9.990000E+2   1.009221E-1   -1.038207E-1   1.300121E-4   -6.770094E-6   6.770094E-6   1.300121E-4   1.301883E-4   -2.980859E+0   8.701914E+1   
9.184110E+2   1.400695E+2   1.400695E+2   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   1.035147E-1   -1.051078E-1   1.324532E-4   -7.846133E-6   7.846133E-6   1.324532E-4   1.326854E-4   -3.390069E+0   8.660993E+1   
9.402480E+2   1.400407E+2   1.400407E+2   8.980000E+2   8.980000E+2   9.000000E+1   8.980000E+2   8.980000E+2   1.039413E-1   -1.060937E-1   1.333591E-4   -7.517102E-6   7.517102E-6   1.333591E-4   1.335708E-4   -3.226199E+0   8.677380E+1   
9.621220E+2   1.398974E+2   1.398974E+2   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   1.040668E-1   -1.075577E-1   1.343901E-4   -6.652796E-6   6.652796E-6   1.343901E-4   1.345547E-4   -2.834034E+0   8.716597E+1   
9.840020E+2   1.400252E+2   1.400252E+2   7.980000E+2   7.980000E+2   9.000000E+1   7.980000E+2   7.980000E+2   1.066648E-1   -1.097317E-1   1.374122E-4   -7.153150E-6   7.153150E-6   1.374122E-4   1.375983E-4   -2.979907E+0   8.702009E+1   
1.005886E+3   1.400380E+2   1.400380E+2   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   1.070568E-1   -1.110116E-1   1.384882E-4   -6.606257E-6   6.606257E-6   1.384882E-4   1.386457E-4   -2.731092E+0   8.726891E+1   
1.027718E+3   1.400487E+2   1.400487E+2   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   1.072555E-1   -1.139499E-1   1.405248E-4   -4.832296E-6   4.832296E-6   1.405248E-4   1.406078E-4   -1.969483E+0   8.803052E+1   
1.049611E+3   1.401052E+2   1.401052E+2   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   1.091653E-1   -1.151726E-1   1.425018E-4   -5.445475E-6   5.445475E-6   1.425018E-4   1.426058E-4   -2.188400E+0   8.781160E+1   
1.071495E+3   1.399861E+2   1.399861E+2   5.980000E+2   5.980000E+2   9.000000E+1   5.990000E+2   5.990000E+2   1.093307E-1   -1.162571E-1   1.433104E-4   -4.858744E-6   4.858744E-6   1.433104E-4   1.433927E-4   -1.941792E+0   8.805821E+1   
1.093324E+3   1.399917E+2   1.399917E+2   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   1.103885E-1   -1.186243E-1   1.455061E-4   -4.093514E-6   4.093514E-6   1.455061E-4   1.455637E-4   -1.611473E+0   8.838853E+1   
1.115201E+3   1.400041E+2   1.400041E+2   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   1.111600E-1   -1.193225E-1   1.464377E-4   -4.207699E-6   4.207699E-6   1.464377E-4   1.464982E-4   -1.645867E+0   8.835413E+1   
1.137095E+3   1.400853E+2   1.400853E+2   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   1.135752E-1   -1.204677E-1   1.486768E-4   -5.245327E-6   5.245327E-6   1.486768E-4   1.487693E-4   -2.020560E+0   8.797944E+1   
1.158972E+3   1.400894E+2   1.400894E+2   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   1.127428E-1   -1.230026E-1   1.498132E-4   -2.972479E-6   2.972479E-6   1.498132E-4   1.498427E-4   -1.136670E+0   8.886333E+1   
1.180841E+3   1.400602E+2   1.400602E+2   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   1.138853E-1   -1.247404E-1   1.516514E-4   -2.681371E-6   2.681371E-6   1.516514E-4   1.516751E-4   -1.012950E+0   8.898705E+1   
1.202710E+3   1.401001E+2   1.401001E+2   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   1.154570E-1   -1.267495E-1   1.539315E-4   -2.530389E-6   2.530389E-6   1.539315E-4   1.539523E-4   -9.417667E-1   8.905823E+1   
1.224513E+3   1.400232E+2   1.400232E+2   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   1.156465E-1   -1.280579E-1   1.549008E-4   -1.815081E-6   1.815081E-6   1.549008E-4   1.549115E-4   -6.713439E-1   8.932866E+1   
1.246394E+3   1.399669E+2   1.399669E+2   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   1.170631E-1   -1.297511E-1   1.568794E-4   -1.755893E-6   1.755893E-6   1.568794E-4   1.568892E-4   -6.412637E-1   8.935874E+1   
1.268274E+3   1.400365E+2   1.400365E+2   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   1.177489E-1   -1.309200E-1   1.580647E-4   -1.498973E-6   1.498973E-6   1.580647E-4   1.580718E-4   -5.433362E-1   8.945666E+1   
1.290111E+3   1.399917E+2   1.399917E+2   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   1.209742E-1   -1.329741E-1   1.613966E-4   -2.541581E-6   2.541581E-6   1.613966E-4   1.614166E-4   -9.021865E-1   8.909781E+1   
1.311842E+3   1.400874E+2   1.400874E+2   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   1.206925E-1   -1.332509E-1   1.614026E-4   -2.152245E-6   2.152245E-6   1.614026E-4   1.614169E-4   -7.639732E-1   8.923603E+1   
1.345031E+3   1.400464E+2   1.400464E+2   4.600000E+1   4.600000E+1   9.000000E+1   4.700000E+1   4.700000E+1   1.190187E-1   -1.335170E-1   1.605412E-4   -7.403141E-7   7.403141E-7   1.605412E-4   1.605429E-4   -2.642100E-1   8.973579E+1   
1.364089E+3   1.400546E+2   1.400546E+2   4.700000E+1   4.700000E+1   9.000000E+1   4.800000E+1   4.800000E+1   1.195041E-1   -1.344038E-1   1.614188E-4   -5.195498E-7   5.195498E-7   1.614188E-4   1.614196E-4   -1.844141E-1   8.981559E+1   
1.386180E+3   1.401434E+2   1.401434E+2   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   1.211467E-1   -1.341734E-1   1.622842E-4   -1.885065E-6   1.885065E-6   1.622842E-4   1.622952E-4   -6.655079E-1   8.933449E+1   
1.405217E+3   1.400603E+2   1.400603E+2   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   1.204835E-1   -1.347538E-1   1.622523E-4   -1.015097E-6   1.015097E-6   1.622523E-4   1.622555E-4   -3.584543E-1   8.964155E+1   
1.427625E+3   1.400797E+2   1.400797E+2   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   1.205311E-1   -1.341376E-1   1.618804E-4   -1.453131E-6   1.453131E-6   1.618804E-4   1.618869E-4   -5.143059E-1   8.948569E+1   
1.446717E+3   1.400128E+2   1.400128E+2   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   1.197978E-1   -1.341395E-1   1.614282E-4   -9.096080E-7   9.096080E-7   1.614282E-4   1.614308E-4   -3.228441E-1   8.967716E+1   
1.469075E+3   1.399924E+2   1.399924E+2   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   1.210887E-1   -1.349016E-1   1.627226E-4   -1.366129E-6   1.366129E-6   1.627226E-4   1.627284E-4   -4.810122E-1   8.951899E+1   
1.488101E+3   1.400740E+2   1.400740E+2   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   1.201663E-1   -1.350063E-1   1.622206E-4   -6.154162E-7   6.154162E-7   1.622206E-4   1.622218E-4   -2.173619E-1   8.978264E+1   
1.510506E+3   1.400219E+2   1.400219E+2   3.100000E+1   3.100000E+1   9.000000E+1   3.100000E+1   3.100000E+1   1.204598E-1   -1.344552E-1   1.620431E-4   -1.192798E-6   1.192798E-6   1.620431E-4   1.620475E-4   -4.217461E-1   8.957825E+1   
1.531906E+3   1.400201E+2   1.400201E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   1.223749E-1   -1.347222E-1   1.634011E-4   -2.434686E-6   2.434686E-6   1.634011E-4   1.634192E-4   -8.536477E-1   8.914635E+1   
1.550969E+3   1.400871E+2   1.400871E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   1.213622E-1   -1.359017E-1   1.635431E-4   -9.145487E-7   9.145487E-7   1.635431E-4   1.635457E-4   -3.204001E-1   8.967960E+1   
1.573411E+3   1.400331E+2   1.400331E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   1.219363E-1   -1.354148E-1   1.635810E-4   -1.657528E-6   1.657528E-6   1.635810E-4   1.635894E-4   -5.805448E-1   8.941946E+1   
1.592440E+3   1.399979E+2   1.399979E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   1.212004E-1   -1.354389E-1   1.631416E-4   -1.097427E-6   1.097427E-6   1.631416E-4   1.631453E-4   -3.854135E-1   8.961459E+1   
1.614867E+3   1.400079E+2   1.400079E+2   2.100000E+1   2.100000E+1   9.000000E+1   2.100000E+1   2.100000E+1   1.234392E-1   -1.353168E-1   1.644463E-4   -2.833158E-6   2.833158E-6   1.644463E-4   1.644707E-4   -9.870213E-1   8.901298E+1   
1.636254E+3   1.400048E+2   1.400048E+2   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   1.222806E-1   -1.353914E-1   1.637785E-4   -1.927464E-6   1.927464E-6   1.637785E-4   1.637899E-4   -6.742669E-1   8.932573E+1   
1.655270E+3   1.400544E+2   1.400544E+2   1.900000E+1   1.900000E+1   9.000000E+1   1.900000E+1   1.900000E+1   1.220108E-1   -1.356027E-1   1.637494E-4   -1.589715E-6   1.589715E-6   1.637494E-4   1.637571E-4   -5.562225E-1   8.944378E+1   
1.677329E+3   1.400093E+2   1.400093E+2   1.500000E+1   1.500000E+1   9.000000E+1   1.500000E+1   1.500000E+1   1.223557E-1   -1.357077E-1   1.640310E-4   -1.776270E-6   1.776270E-6   1.640310E-4   1.640406E-4   -6.204242E-1   8.937958E+1   
1.698740E+3   1.400002E+2   1.400002E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   1.221456E-1   -1.356438E-1   1.638595E-4   -1.662564E-6   1.662564E-6   1.638595E-4   1.638679E-4   -5.813190E-1   8.941868E+1   
1.717838E+3   1.400669E+2   1.400669E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   1.213988E-1   -1.363130E-1   1.638336E-4   -6.728032E-7   6.728032E-7   1.638336E-4   1.638350E-4   -2.352909E-1   8.976471E+1   
1.739931E+3   1.400418E+2   1.400418E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   1.228360E-1   -1.350258E-1   1.638838E-4   -2.577280E-6   2.577280E-6   1.638838E-4   1.639041E-4   -9.009740E-1   8.909903E+1   
1.758597E+3   1.401334E+2   1.401334E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   1.218162E-1   -1.355934E-1   1.636230E-4   -1.451961E-6   1.451961E-6   1.636230E-4   1.636295E-4   -5.084190E-1   8.949158E+1   
1.780579E+3   1.399851E+2   1.399851E+2   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   1.214129E-1   -1.371529E-1   1.643894E-4   -1.340667E-7   1.340667E-7   1.643894E-4   1.643895E-4   -4.672719E-2   8.995327E+1   
1.799249E+3   1.400153E+2   1.400153E+2   5.000000E+0   5.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   1.227702E-1   -1.357800E-1   1.643344E-4   -2.035499E-6   2.035499E-6   1.643344E-4   1.643470E-4   -7.096480E-1   8.929035E+1   
1.820978E+3   1.400164E+2   1.400164E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   1.215740E-1   -1.374150E-1   1.646596E-4   -8.190928E-8   8.190928E-8   1.646596E-4   1.646597E-4   -2.850155E-2   8.997150E+1   
1.839742E+3   1.400470E+2   1.400470E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   1.223203E-1   -1.364855E-1   1.645157E-4   -1.241513E-6   1.241513E-6   1.645157E-4   1.645204E-4   -4.323728E-1   8.956763E+1   
1.861730E+3   1.400037E+2   1.400037E+2   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   1.232695E-1   -1.359345E-1   1.647437E-4   -2.303812E-6   2.303812E-6   1.647437E-4   1.647598E-4   -8.011846E-1   8.919882E+1   
1.883746E+3   1.400381E+2   1.400381E+2   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   1.235060E-1   -1.360031E-1   1.649346E-4   -2.433917E-6   2.433917E-6   1.649346E-4   1.649525E-4   -8.454446E-1   8.915456E+1   
1.905844E+3   1.400488E+2   1.400488E+2   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   1.229268E-1   -1.368178E-1   1.651071E-4   -1.472901E-6   1.472901E-6   1.651071E-4   1.651137E-4   -5.111154E-1   8.948888E+1   
1.927839E+3   1.400141E+2   1.400141E+2   -8.000000E+0   -8.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   1.230434E-1   -1.362797E-1   1.648287E-4   -1.910922E-6   1.910922E-6   1.648287E-4   1.648398E-4   -6.642221E-1   8.933578E+1   
1.949896E+3   1.400679E+2   1.400679E+2   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   1.229121E-1   -1.377133E-1   1.656812E-4   -8.765416E-7   8.765416E-7   1.656812E-4   1.656835E-4   -3.031222E-1   8.969688E+1   
1.972158E+3   1.400153E+2   1.400153E+2   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   1.238618E-1   -1.371638E-1   1.659105E-4   -1.938175E-6   1.938175E-6   1.659105E-4   1.659218E-4   -6.693019E-1   8.933070E+1   
1.994439E+3   1.400337E+2   1.400337E+2   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   1.227658E-1   -1.370235E-1   1.651415E-4   -1.219291E-6   1.219291E-6   1.651415E-4   1.651460E-4   -4.230250E-1   8.957698E+1   
2.016671E+3   1.400224E+2   1.400224E+2   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   1.233881E-1   -1.370287E-1   1.655296E-4   -1.676167E-6   1.676167E-6   1.655296E-4   1.655381E-4   -5.801620E-1   8.941984E+1   
2.038934E+3   1.400926E+2   1.400926E+2   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   1.246791E-1   -1.364398E-1   1.659442E-4   -3.016021E-6   3.016021E-6   1.659442E-4   1.659716E-4   -1.041231E+0   8.895877E+1   
2.061200E+3   1.399770E+2   1.399770E+2   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   1.228675E-1   -1.361573E-1   1.646402E-4   -1.860814E-6   1.860814E-6   1.646402E-4   1.646507E-4   -6.475470E-1   8.935245E+1   
2.083467E+3   1.399972E+2   1.399972E+2   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   1.228843E-1   -1.368441E-1   1.650980E-4   -1.424238E-6   1.424238E-6   1.650980E-4   1.651041E-4   -4.942568E-1   8.950574E+1   
2.105713E+3   1.399826E+2   1.399826E+2   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   1.239757E-1   -1.375323E-1   1.662209E-4   -1.781577E-6   1.781577E-6   1.662209E-4   1.662305E-4   -6.140799E-1   8.938592E+1   
2.127962E+3   1.400585E+2   1.400585E+2   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   1.236199E-1   -1.384293E-1   1.665852E-4   -9.319071E-7   9.319071E-7   1.665852E-4   1.665878E-4   -3.205195E-1   8.967948E+1   
2.150232E+3   1.400769E+2   1.400769E+2   -2.700000E+1   -2.700000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   1.241796E-1   -1.382322E-1   1.668028E-4   -1.474764E-6   1.474764E-6   1.668028E-4   1.668094E-4   -5.065593E-1   8.949344E+1   
2.172144E+3   1.399735E+2   1.399735E+2   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   1.228972E-1   -1.376328E-1   1.656196E-4   -9.181856E-7   9.181856E-7   1.656196E-4   1.656221E-4   -3.176413E-1   8.968236E+1   
2.194337E+3   1.400858E+2   1.400858E+2   -3.100000E+1   -3.100000E+1   9.000000E+1   -3.000000E+1   -3.000000E+1   1.247297E-1   -1.380712E-1   1.670380E-4   -1.986914E-6   1.986914E-6   1.670380E-4   1.670498E-4   -6.815001E-1   8.931850E+1   
2.216259E+3   1.399444E+2   1.399444E+2   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   1.238587E-1   -1.381962E-1   1.665810E-4   -1.260969E-6   1.260969E-6   1.665810E-4   1.665857E-4   -4.337041E-1   8.956630E+1   
2.238479E+3   1.400219E+2   1.400219E+2   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   1.241729E-1   -1.384148E-1   1.669176E-4   -1.350431E-6   1.350431E-6   1.669176E-4   1.669230E-4   -4.635359E-1   8.953646E+1   
2.260746E+3   1.399650E+2   1.399650E+2   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   1.228926E-1   -1.392522E-1   1.666714E-4   1.439443E-7   -1.439443E-7   1.666714E-4   1.666715E-4   4.948297E-2   9.004948E+1   
2.283040E+3   1.400527E+2   1.400527E+2   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   1.234432E-1   -1.388119E-1   1.667251E-4   -5.510892E-7   5.510892E-7   1.667251E-4   1.667260E-4   -1.893834E-1   8.981062E+1   
2.305285E+3   1.400641E+2   1.400641E+2   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   1.237658E-1   -1.386252E-1   1.668029E-4   -9.117341E-7   9.117341E-7   1.668029E-4   1.668054E-4   -3.131719E-1   8.968683E+1   
2.327523E+3   1.400595E+2   1.400595E+2   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   1.246610E-1   -1.384939E-1   1.672709E-4   -1.659699E-6   1.659699E-6   1.672709E-4   1.672791E-4   -5.684829E-1   8.943152E+1   
2.349767E+3   1.399929E+2   1.399929E+2   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   1.249587E-1   -1.385077E-1   1.674639E-4   -1.870898E-6   1.870898E-6   1.674639E-4   1.674744E-4   -6.400785E-1   8.935992E+1   
2.372039E+3   1.399727E+2   1.399727E+2   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   1.238983E-1   -1.392325E-1   1.672804E-4   -6.127238E-7   6.127238E-7   1.672804E-4   1.672815E-4   -2.098652E-1   8.979013E+1   
2.394311E+3   1.400059E+2   1.400059E+2   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   1.257096E-1   -1.384297E-1   1.678773E-4   -2.477317E-6   2.477317E-6   1.678773E-4   1.678956E-4   -8.454360E-1   8.915456E+1   
2.427674E+3   1.401072E+2   1.401072E+2   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   1.264287E-1   -1.403447E-1   1.695691E-4   -1.757212E-6   1.757212E-6   1.695691E-4   1.695782E-4   -5.937238E-1   8.940628E+1   
2.449389E+3   1.400368E+2   1.400368E+2   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   1.261316E-1   -1.434640E-1   1.714170E-4   5.018710E-7   -5.018710E-7   1.714170E-4   1.714177E-4   1.677489E-1   9.016775E+1   
2.471079E+3   1.399786E+2   1.399786E+2   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   1.283498E-1   -1.434641E-1   1.727885E-4   -1.138739E-6   1.138739E-6   1.727885E-4   1.727923E-4   -3.775943E-1   8.962241E+1   
2.492744E+3   1.400225E+2   1.400225E+2   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   1.292627E-1   -1.445259E-1   1.740445E-4   -1.119732E-6   1.119732E-6   1.740445E-4   1.740481E-4   -3.686128E-1   8.963139E+1   
2.514437E+3   1.399744E+2   1.399744E+2   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   1.305228E-1   -1.461306E-1   1.758687E-4   -1.002683E-6   1.002683E-6   1.758687E-4   1.758715E-4   -3.266580E-1   8.967334E+1   
2.536120E+3   1.399793E+2   1.399793E+2   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   1.309524E-1   -1.472688E-1   1.768755E-4   -5.762510E-7   5.762510E-7   1.768755E-4   1.768764E-4   -1.866660E-1   8.981333E+1   
2.557807E+3   1.399391E+2   1.399391E+2   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   1.314641E-1   -1.500076E-1   1.789756E-4   8.357797E-7   -8.357797E-7   1.789756E-4   1.789775E-4   2.675577E-1   9.026756E+1   
2.580049E+3   1.400133E+2   1.400133E+2   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   1.328014E-1   -1.505610E-1   1.801628E-4   2.084880E-7   -2.084880E-7   1.801628E-4   1.801629E-4   6.630380E-2   9.006630E+1   
2.601736E+3   1.400316E+2   1.400316E+2   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   1.330994E-1   -1.524205E-1   1.815581E-4   1.203728E-6   -1.203728E-6   1.815581E-4   1.815621E-4   3.798645E-1   9.037986E+1   
2.623465E+3   1.400904E+2   1.400904E+2   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   1.347675E-1   -1.534364E-1   1.832511E-4   6.341713E-7   -6.341713E-7   1.832511E-4   1.832522E-4   1.982810E-1   9.019828E+1   
2.645142E+3   1.401270E+2   1.401270E+2   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   1.350125E-1   -1.546441E-1   1.841891E-4   1.242543E-6   -1.242543E-6   1.841891E-4   1.841933E-4   3.865125E-1   9.038651E+1   
2.666889E+3   1.400184E+2   1.400184E+2   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.500000E+2   -6.500000E+2   1.348222E-1   -1.558220E-1   1.848386E-4   2.153332E-6   -2.153332E-6   1.848386E-4   1.848512E-4   6.674537E-1   9.066745E+1   
2.688606E+3   1.400747E+2   1.400747E+2   -7.000000E+2   -7.000000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   1.374608E-1   -1.587672E-1   1.883881E-4   2.127262E-6   -2.127262E-6   1.883881E-4   1.884001E-4   6.469514E-1   9.064695E+1   
2.710347E+3   1.400063E+2   1.400063E+2   -7.510000E+2   -7.510000E+2   9.000000E+1   -7.490000E+2   -7.490000E+2   1.373401E-1   -1.599935E-1   1.891121E-4   3.018226E-6   -3.018226E-6   1.891121E-4   1.891362E-4   9.143619E-1   9.091436E+1   
2.732077E+3   1.400395E+2   1.400395E+2   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   1.388828E-1   -1.611544E-1   1.908220E-4   2.636170E-6   -2.636170E-6   1.908220E-4   1.908402E-4   7.914800E-1   9.079148E+1   
2.753804E+3   1.399710E+2   1.399710E+2   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   1.388641E-1   -1.634724E-1   1.923201E-4   4.165421E-6   -4.165421E-6   1.923201E-4   1.923652E-4   1.240764E+0   9.124076E+1   
2.775508E+3   1.400061E+2   1.400061E+2   -9.000000E+2   -9.000000E+2   9.000000E+1   -9.000000E+2   -9.000000E+2   1.402457E-1   -1.654981E-1   1.944936E-4   4.467899E-6   -4.467899E-6   1.944936E-4   1.945449E-4   1.315965E+0   9.131596E+1   
2.797242E+3   1.400151E+2   1.400151E+2   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.490000E+2   -9.490000E+2   1.404349E-1   -1.669586E-1   1.955618E-4   5.282838E-6   -5.282838E-6   1.955618E-4   1.956331E-4   1.547392E+0   9.154739E+1   
2.818977E+3   1.400313E+2   1.400313E+2   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   1.428670E-1   -1.683611E-1   1.979789E-4   4.400902E-6   -4.400902E-6   1.979789E-4   1.980278E-4   1.273427E+0   9.127343E+1   
2.841096E+3   1.400296E+2   1.400296E+2   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   1.436632E-1   -1.687394E-1   1.987175E-4   4.059260E-6   -4.059260E-6   1.987175E-4   1.987590E-4   1.170235E+0   9.117023E+1   
2.862868E+3   1.400256E+2   1.400256E+2   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   1.444258E-1   -1.706266E-1   2.004181E-4   4.729085E-6   -4.729085E-6   2.004181E-4   2.004739E-4   1.351706E+0   9.135171E+1   
2.884685E+3   1.399566E+2   1.399566E+2   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   1.463125E-1   -1.719759E-1   2.024633E-4   4.215691E-6   -4.215691E-6   2.024633E-4   2.025072E-4   1.192840E+0   9.119284E+1   
2.907208E+3   1.400803E+2   1.400803E+2   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   1.464725E-1   -1.746505E-1   2.043042E-4   5.845928E-6   -5.845928E-6   2.043042E-4   2.043878E-4   1.639005E+0   9.163900E+1   
2.929285E+3   1.400695E+2   1.400695E+2   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   1.472608E-1   -1.759943E-1   2.056667E-4   6.141390E-6   -6.141390E-6   2.056667E-4   2.057584E-4   1.710394E+0   9.171039E+1   
2.951407E+3   1.399907E+2   1.399907E+2   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   1.480613E-1   -1.765689E-1   2.065358E-4   5.925044E-6   -5.925044E-6   2.065358E-4   2.066208E-4   1.643235E+0   9.164324E+1   
2.974021E+3   1.400502E+2   1.400502E+2   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   1.482137E-1   -1.788987E-1   2.081474E-4   7.335419E-6   -7.335419E-6   2.081474E-4   2.082767E-4   2.018351E+0   9.201835E+1   
2.996143E+3   1.400012E+2   1.400012E+2   -1.399000E+3   -1.399000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   1.490275E-1   -1.802443E-1   2.095269E-4   7.613232E-6   -7.613232E-6   2.095269E-4   2.096652E-4   2.080946E+0   9.208095E+1   
3.018278E+3   1.400371E+2   1.400371E+2   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   1.502872E-1   -1.814078E-1   2.110635E-4   7.442212E-6   -7.442212E-6   2.110635E-4   2.111947E-4   2.019443E+0   9.201944E+1   
3.040661E+3   1.399834E+2   1.399834E+2   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   1.529808E-1   -1.829044E-1   2.137036E-4   6.428321E-6   -6.428321E-6   2.137036E-4   2.138002E-4   1.722969E+0   9.172297E+1   
3.062779E+3   1.400798E+2   1.400798E+2   -1.550000E+3   -1.550000E+3   9.000000E+1   -1.548000E+3   -1.548000E+3   1.520230E-1   -1.848290E-1   2.143649E-4   8.395004E-6   -8.395004E-6   2.143649E-4   2.145292E-4   2.242683E+0   9.224268E+1   
3.084941E+3   1.400560E+2   1.400560E+2   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   1.538156E-1   -1.855456E-1   2.159399E-4   7.537648E-6   -7.537648E-6   2.159399E-4   2.160714E-4   1.999168E+0   9.199917E+1   
3.107790E+3   1.400453E+2   1.400453E+2   -1.650000E+3   -1.650000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   1.551560E-1   -1.881967E-1   2.184952E-4   8.279525E-6   -8.279525E-6   2.184952E-4   2.186521E-4   2.170093E+0   9.217009E+1   
3.129860E+3   1.399891E+2   1.399891E+2   -1.700000E+3   -1.700000E+3   9.000000E+1   -1.698000E+3   -1.698000E+3   1.557844E-1   -1.886356E-1   2.191696E-4   8.101584E-6   -8.101584E-6   2.191696E-4   2.193193E-4   2.116970E+0   9.211697E+1   
3.151901E+3   1.400319E+2   1.400319E+2   -1.750000E+3   -1.750000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   1.579740E-1   -1.907108E-1   2.218748E-4   7.838807E-6   -7.838807E-6   2.218748E-4   2.220133E-4   2.023410E+0   9.202341E+1   
3.174945E+3   1.399864E+2   1.399864E+2   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.799000E+3   -1.799000E+3   1.580941E-1   -1.919879E-1   2.227809E-4   8.584931E-6   -8.584931E-6   2.227809E-4   2.229462E-4   2.206819E+0   9.220682E+1   
3.197018E+3   1.399921E+2   1.399921E+2   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.848000E+3   -1.848000E+3   1.591365E-1   -1.940628E-1   2.247766E-4   9.170473E-6   -9.170473E-6   2.247766E-4   2.249636E-4   2.336267E+0   9.233627E+1   
3.219088E+3   1.399751E+2   1.399751E+2   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   1.610107E-1   -1.961991E-1   2.273267E-4   9.180950E-6   -9.180950E-6   2.273267E-4   2.275121E-4   2.312724E+0   9.231272E+1   
3.242370E+3   1.400709E+2   1.400709E+2   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.948000E+3   -1.948000E+3   1.606974E-1   -1.973079E-1   2.278552E-4   1.013749E-5   -1.013749E-5   2.278552E-4   2.280806E-4   2.547462E+0   9.254746E+1   
3.264491E+3   1.399900E+2   1.399900E+2   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   1.626799E-1   -2.001966E-1   2.309623E-4   1.055978E-5   -1.055978E-5   2.309623E-4   2.312036E-4   2.617786E+0   9.261779E+1   
3.301612E+3   1.400603E+2   1.400603E+2   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.711023E-1   -2.149343E-1   2.457679E-4   1.396541E-5   -1.396541E-5   2.457679E-4   2.461644E-4   3.252254E+0   9.325225E+1   
3.327734E+3   1.400260E+2   1.400260E+2   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.800489E-1   -2.302425E-1   2.612691E-4   1.735633E-5   -1.735633E-5   2.612691E-4   2.618450E-4   3.800623E+0   9.380062E+1   
3.353900E+3   1.400200E+2   1.400200E+2   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.906687E-1   -2.460960E-1   2.781600E-4   1.986613E-5   -1.986613E-5   2.781600E-4   2.788685E-4   4.085117E+0   9.408512E+1   
3.379600E+3   1.399986E+2   1.399986E+2   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   1.941996E-1   -2.552660E-1   2.863153E-4   2.324965E-5   -2.324965E-5   2.863153E-4   2.872577E-4   4.642401E+0   9.464240E+1   
3.405341E+3   1.400258E+2   1.400258E+2   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   1.926800E-1   -2.594909E-1   2.881274E-4   2.713573E-5   -2.713573E-5   2.881274E-4   2.894024E-4   5.380225E+0   9.538022E+1   
3.430088E+3   1.400051E+2   1.400051E+2   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   1.775416E-1   -2.467878E-1   2.704947E-4   3.002762E-5   -3.002762E-5   2.704947E-4   2.721563E-4   6.334469E+0   9.633447E+1   
3.455347E+3   1.399568E+2   1.399568E+2   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   1.599314E-1   -2.279946E-1   2.473675E-4   3.076624E-5   -3.076624E-5   2.473675E-4   2.492735E-4   7.089731E+0   9.708973E+1   
3.481043E+3   1.399889E+2   1.399889E+2   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   1.447602E-1   -2.128786E-1   2.281431E-4   3.210492E-5   -3.210492E-5   2.281431E-4   2.303910E-4   8.010219E+0   9.801022E+1   
3.505794E+3   1.399301E+2   1.399301E+2   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.363949E-1   -2.078675E-1   2.197076E-4   3.501603E-5   -3.501603E-5   2.197076E-4   2.224804E-4   9.055392E+0   9.905539E+1   
3.530536E+3   1.400505E+2   1.400505E+2   -7.001000E+3   -7.001000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.327566E-1   -2.044109E-1   2.152070E-4   3.544714E-5   -3.544714E-5   2.152070E-4   2.181067E-4   9.353314E+0   9.935331E+1   
3.555739E+3   1.400442E+2   1.400442E+2   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.360924E-1   -2.139936E-1   2.235104E-4   3.924480E-5   -3.924480E-5   2.235104E-4   2.269296E-4   9.958695E+0   9.995870E+1   
3.580939E+3   1.400470E+2   1.400470E+2   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.380905E-1   -2.209157E-1   2.292541E-4   4.229243E-5   -4.229243E-5   2.292541E-4   2.331224E-4   1.045232E+1   1.004523E+2   
3.606162E+3   1.400117E+2   1.400117E+2   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.500000E+3   -8.500000E+3   1.456379E-1   -2.348432E-1   2.429910E-4   4.581552E-5   -4.581552E-5   2.429910E-4   2.472725E-4   1.067766E+1   1.006777E+2   
3.631872E+3   1.400591E+2   1.400591E+2   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.633555E-1   -2.566805E-1   2.681673E-4   4.698769E-5   -4.698769E-5   2.681673E-4   2.722527E-4   9.938354E+0   9.993835E+1   
3.657105E+3   1.400568E+2   1.400568E+2   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.732606E-1   -2.706882E-1   2.834142E-4   4.881942E-5   -4.881942E-5   2.834142E-4   2.875881E-4   9.773554E+0   9.977355E+1   
3.682352E+3   1.399582E+2   1.399582E+2   -9.999000E+3   -9.999000E+3   9.000000E+1   -9.999000E+3   -9.999000E+3   1.834719E-1   -2.890485E-1   3.016852E-4   5.327021E-5   -5.327021E-5   3.016852E-4   3.063522E-4   1.001381E+1   1.000138E+2   
3.718887E+3   1.400060E+2   1.400060E+2   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.731093E-1   -2.698144E-1   2.827515E-4   4.836000E-5   -4.836000E-5   2.827515E-4   2.868573E-4   9.705590E+0   9.970559E+1   
3.743062E+3   1.399803E+2   1.399803E+2   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.566312E-1   -2.496461E-1   2.594286E-4   4.736225E-5   -4.736225E-5   2.594286E-4   2.637165E-4   1.034619E+1   1.003462E+2   
3.767797E+3   1.399519E+2   1.399519E+2   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.454287E-1   -2.325177E-1   2.413471E-4   4.444994E-5   -4.444994E-5   2.413471E-4   2.454062E-4   1.043547E+1   1.004355E+2   
3.792471E+3   1.399905E+2   1.399905E+2   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.383835E-1   -2.190808E-1   2.282401E-4   4.087611E-5   -4.087611E-5   2.282401E-4   2.318715E-4   1.015360E+1   1.001536E+2   
3.817240E+3   1.400251E+2   1.400251E+2   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.258728E-1   -2.010678E-1   2.087737E-4   3.835298E-5   -3.835298E-5   2.087737E-4   2.122674E-4   1.040951E+1   1.004095E+2   
3.842337E+3   1.400946E+2   1.400946E+2   -7.000000E+3   -7.000000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.146825E-1   -1.829522E-1   1.900569E-4   3.478621E-5   -3.478621E-5   1.900569E-4   1.932142E-4   1.037207E+1   1.003721E+2   
3.867075E+3   1.400454E+2   1.400454E+2   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.049241E-1   -1.661494E-1   1.730803E-4   3.101871E-5   -3.101871E-5   1.730803E-4   1.758379E-4   1.016044E+1   1.001604E+2   
3.891284E+3   1.399601E+2   1.399601E+2   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   9.271197E-2   -1.492237E-1   1.545067E-4   2.898559E-5   -2.898559E-5   1.545067E-4   1.572020E-4   1.062524E+1   1.006252E+2   
3.916025E+3   1.399811E+2   1.399811E+2   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   8.235574E-2   -1.310827E-1   1.362890E-4   2.478533E-5   -2.478533E-5   1.362890E-4   1.385244E-4   1.030709E+1   1.003071E+2   
3.941172E+3   1.400693E+2   1.400693E+2   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   7.140601E-2   -1.144813E-1   1.187070E-4   2.203053E-5   -2.203053E-5   1.187070E-4   1.207340E-4   1.051376E+1   1.005138E+2   
3.965918E+3   1.400266E+2   1.400266E+2   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   5.978501E-2   -9.746468E-2   1.004396E-4   1.950080E-5   -1.950080E-5   1.004396E-4   1.023152E-4   1.098753E+1   1.009875E+2   
3.990512E+3   1.400286E+2   1.400286E+2   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   4.879691E-2   -8.158172E-2   8.330184E-5   1.724411E-5   -1.724411E-5   8.330184E-5   8.506795E-5   1.169547E+1   1.016955E+2   
4.015224E+3   1.399640E+2   1.399640E+2   -3.499000E+3   -3.499000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   3.809125E-2   -6.178900E-2   6.379231E-5   1.222243E-5   -1.222243E-5   6.379231E-5   6.495265E-5   1.084627E+1   1.008463E+2   
4.039417E+3   1.400546E+2   1.400546E+2   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   2.696047E-2   -4.581543E-2   4.650732E-5   1.001203E-5   -1.001203E-5   4.650732E-5   4.757281E-5   1.214914E+1   1.021491E+2   
4.064602E+3   1.399748E+2   1.399748E+2   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.658407E-2   -2.986456E-2   2.970352E-5   7.258517E-6   -7.258517E-6   2.970352E-5   3.057753E-5   1.373200E+1   1.037320E+2   
4.089294E+3   1.400330E+2   1.400330E+2   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   7.930016E-3   -1.265036E-2   1.314175E-5   2.405163E-6   -2.405163E-6   1.314175E-5   1.336003E-5   1.037132E+1   1.003713E+2   
4.122955E+3   1.400406E+2   1.400406E+2   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   6.084035E-3   -9.348020E-3   9.849701E-6   1.611530E-6   -1.611530E-6   9.849701E-6   9.980663E-6   9.291953E+0   9.929195E+1   
4.145047E+3   1.400111E+2   1.400111E+2   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   3.954576E-3   -8.870951E-3   8.222460E-6   2.874650E-6   -2.874650E-6   8.222460E-6   8.710480E-6   1.927011E+1   1.092701E+2   
4.167083E+3   1.400526E+2   1.400526E+2   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.849000E+3   -1.849000E+3   4.060115E-3   -6.159814E-3   6.521975E-6   1.024126E-6   -1.024126E-6   6.521975E-6   6.601893E-6   8.924108E+0   9.892411E+1   
4.188868E+3   1.400732E+2   1.400732E+2   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.799000E+3   -1.799000E+3   2.749795E-3   -3.799647E-3   4.174722E-6   4.502678E-7   -4.502678E-7   4.174722E-6   4.198934E-6   6.155883E+0   9.615588E+1   
4.210863E+3   1.400040E+2   1.400040E+2   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   3.874804E-4   -4.050910E-3   2.877873E-6   2.361778E-6   -2.361778E-6   2.877873E-6   3.722922E-6   3.937463E+1   1.293746E+2   
4.232861E+3   1.401121E+2   1.401121E+2   -1.700000E+3   -1.700000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   4.835088E-4   -1.097403E-3   1.013655E-6   3.598332E-7   -3.598332E-7   1.013655E-6   1.075628E-6   1.954414E+1   1.095441E+2   
4.254657E+3   1.400963E+2   1.400963E+2   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   -6.227917E-4   -1.733385E-4   -2.721454E-7   5.739599E-7   -5.739599E-7   -2.721454E-7   6.352111E-7   1.153682E+2   2.053682E+2   
4.276477E+3   1.400425E+2   1.400425E+2   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   -2.705926E-3   1.881569E-3   -2.898376E-6   7.712703E-7   -7.712703E-7   -2.898376E-6   2.999240E-6   1.650987E+2   2.550987E+2   
4.298345E+3   1.401534E+2   1.401534E+2   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   -2.667883E-3   4.272724E-3   -4.432190E-6   -8.201374E-7   8.201374E-7   -4.432190E-6   4.507431E-6   -1.695165E+2   -7.951650E+1   
4.320185E+3   1.400542E+2   1.400542E+2   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   -3.211524E-3   5.632743E-3   -5.654060E-6   -1.307186E-6   1.307186E-6   -5.654060E-6   5.803200E-6   -1.669823E+2   -7.698227E+1   
4.342299E+3   1.400011E+2   1.400011E+2   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   -5.653604E-3   7.998123E-3   -8.704415E-6   -1.047366E-6   1.047366E-6   -8.704415E-6   8.767201E-6   -1.731388E+2   -8.313882E+1   
4.364399E+3   1.400350E+2   1.400350E+2   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   -5.859769E-3   8.954400E-3   -9.454689E-6   -1.520067E-6   1.520067E-6   -9.454689E-6   9.576103E-6   -1.708665E+2   -8.086650E+1   
4.386173E+3   1.399853E+2   1.399853E+2   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.350000E+3   -1.350000E+3   -7.103820E-3   1.078014E-2   -1.141290E-5   -1.793542E-6   1.793542E-6   -1.141290E-5   1.155297E-5   -1.710690E+2   -8.106899E+1   
4.408228E+3   1.399473E+2   1.399473E+2   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   -8.116547E-3   1.120474E-2   -1.231556E-5   -1.322093E-6   1.322093E-6   -1.231556E-5   1.238632E-5   -1.738727E+2   -8.387268E+1   
4.430293E+3   1.400429E+2   1.400429E+2   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.250000E+3   -1.250000E+3   -7.641018E-3   1.458009E-2   -1.421990E-5   -3.880519E-6   3.880519E-6   -1.421990E-5   1.473987E-5   -1.647360E+2   -7.473601E+1   
4.452365E+3   1.399549E+2   1.399549E+2   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   -1.025214E-2   1.592876E-2   -1.671259E-5   -2.830970E-6   2.830970E-6   -1.671259E-5   1.695066E-5   -1.703858E+2   -8.038584E+1   
4.474452E+3   1.399879E+2   1.399879E+2   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.150000E+3   -1.150000E+3   -1.108662E-2   1.751641E-2   -1.826252E-5   -3.251727E-6   3.251727E-6   -1.826252E-5   1.854976E-5   -1.699040E+2   -7.990403E+1   
4.496481E+3   1.399832E+2   1.399832E+2   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.100000E+3   -1.100000E+3   -1.146214E-2   1.855184E-2   -1.916905E-5   -3.650911E-6   3.650911E-6   -1.916905E-5   1.951362E-5   -1.692167E+2   -7.921667E+1   
4.518470E+3   1.400398E+2   1.400398E+2   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.050000E+3   -1.050000E+3   -1.182385E-2   2.009285E-2   -2.039632E-5   -4.390851E-6   4.390851E-6   -2.039632E-5   2.086359E-5   -1.678510E+2   -7.785097E+1   
4.540494E+3   1.400169E+2   1.400169E+2   -1.000000E+3   -1.000000E+3   9.000000E+1   -1.000000E+3   -1.000000E+3   -1.423802E-2   2.107583E-2   -2.252907E-5   -3.247905E-6   3.247905E-6   -2.252907E-5   2.276199E-5   -1.717965E+2   -8.179647E+1   
4.562376E+3   1.400708E+2   1.400708E+2   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   -1.541979E-2   2.352591E-2   -2.485541E-5   -3.975624E-6   3.975624E-6   -2.485541E-5   2.517136E-5   -1.709125E+2   -8.091252E+1   
4.583992E+3   1.400782E+2   1.400782E+2   -9.000000E+2   -9.000000E+2   9.000000E+1   -9.000000E+2   -9.000000E+2   -1.632974E-2   2.531393E-2   -2.658250E-5   -4.471549E-6   4.471549E-6   -2.658250E-5   2.695596E-5   -1.704514E+2   -8.045144E+1   
4.605871E+3   1.400695E+2   1.400695E+2   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   -1.662824E-2   2.608429E-2   -2.726878E-5   -4.754405E-6   4.754405E-6   -2.726878E-5   2.768015E-5   -1.701097E+2   -8.010970E+1   
4.627483E+3   1.399384E+2   1.399384E+2   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   -1.810576E-2   2.752930E-2   -2.912337E-5   -4.606296E-6   4.606296E-6   -2.912337E-5   2.948540E-5   -1.710123E+2   -8.101227E+1   
4.649111E+3   1.400483E+2   1.400483E+2   -7.510000E+2   -7.510000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   -1.947835E-2   2.998363E-2   -3.157045E-5   -5.195654E-6   5.195654E-6   -3.157045E-5   3.199513E-5   -1.706544E+2   -8.065441E+1   
4.671046E+3   1.400277E+2   1.400277E+2   -7.000000E+2   -7.000000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   -1.961550E-2   3.067607E-2   -3.210622E-5   -5.546914E-6   5.546914E-6   -3.210622E-5   3.258186E-5   -1.701979E+2   -8.019791E+1   
4.692979E+3   1.400265E+2   1.400265E+2   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.500000E+2   -6.500000E+2   -2.004624E-2   3.300830E-2   -3.389148E-5   -6.753076E-6   6.753076E-6   -3.389148E-5   3.455773E-5   -1.687311E+2   -7.873107E+1   
4.714667E+3   1.401179E+2   1.401179E+2   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   -2.272056E-2   3.474046E-2   -3.667301E-5   -5.907498E-6   5.907498E-6   -3.667301E-5   3.714577E-5   -1.708491E+2   -8.084908E+1   
4.736291E+3   1.400386E+2   1.400386E+2   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   -2.267393E-2   3.634499E-2   -3.768919E-5   -6.990983E-6   6.990983E-6   -3.768919E-5   3.833209E-5   -1.694916E+2   -7.949162E+1   
4.757955E+3   1.399983E+2   1.399983E+2   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   -2.337741E-2   3.703280E-2   -3.857208E-5   -6.920339E-6   6.920339E-6   -3.857208E-5   3.918796E-5   -1.698286E+2   -7.982860E+1   
4.779629E+3   1.400899E+2   1.400899E+2   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   -2.527127E-2   3.849223E-2   -4.069346E-5   -6.473714E-6   6.473714E-6   -4.069346E-5   4.120518E-5   -1.709609E+2   -8.096086E+1   
4.801257E+3   1.400624E+2   1.400624E+2   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   -2.469819E-2   3.951445E-2   -4.100492E-5   -7.565882E-6   7.565882E-6   -4.100492E-5   4.169707E-5   -1.695458E+2   -7.954584E+1   
4.822931E+3   1.400884E+2   1.400884E+2   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   -2.629076E-2   4.229860E-2   -4.380280E-5   -8.208164E-6   8.208164E-6   -4.380280E-5   4.456523E-5   -1.693865E+2   -7.938649E+1   
4.844563E+3   1.399694E+2   1.399694E+2   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   -2.722955E-2   4.308306E-2   -4.489412E-5   -8.026668E-6   8.026668E-6   -4.489412E-5   4.560602E-5   -1.698631E+2   -7.986313E+1   
4.866207E+3   1.399915E+2   1.399915E+2   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   -2.856992E-2   4.471921E-2   -4.678841E-5   -8.104955E-6   8.104955E-6   -4.678841E-5   4.748521E-5   -1.701724E+2   -8.017242E+1   
4.887829E+3   1.400467E+2   1.400467E+2   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   -2.881965E-2   4.703219E-2   -4.844922E-5   -9.432413E-6   9.432413E-6   -4.844922E-5   4.935886E-5   -1.689831E+2   -7.898309E+1   
4.909431E+3   1.400056E+2   1.400056E+2   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   -2.974586E-2   4.699168E-2   -4.899546E-5   -8.720876E-6   8.720876E-6   -4.899546E-5   4.976554E-5   -1.699074E+2   -7.990742E+1   
4.931118E+3   1.401026E+2   1.401026E+2   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   -3.085063E-2   4.960224E-2   -5.137872E-5   -9.610460E-6   9.610460E-6   -5.137872E-5   5.226982E-5   -1.694052E+2   -7.940518E+1   
4.952690E+3   1.400197E+2   1.400197E+2   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   -3.259534E-2   5.021397E-2   -5.285580E-5   -8.719949E-6   8.719949E-6   -5.285580E-5   5.357026E-5   -1.706319E+2   -8.063194E+1   
4.985731E+3   1.400257E+2   1.400257E+2   -4.700000E+1   -4.700000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   -3.204590E-2   5.111567E-2   -5.310337E-5   -9.715838E-6   9.715838E-6   -5.310337E-5   5.398486E-5   -1.696318E+2   -7.963179E+1   
5.007018E+3   1.400382E+2   1.400382E+2   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   -3.215141E-2   5.122551E-2   -5.324014E-5   -9.709609E-6   9.709609E-6   -5.324014E-5   5.411829E-5   -1.696643E+2   -7.966434E+1   
5.029210E+3   1.400400E+2   1.400400E+2   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   -3.251345E-2   5.023916E-2   -5.282157E-5   -8.796986E-6   8.796986E-6   -5.282157E-5   5.354910E-5   -1.705447E+2   -8.054465E+1   
5.051448E+3   1.400243E+2   1.400243E+2   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   -3.190046E-2   5.138535E-2   -5.318909E-5   -9.999715E-6   9.999715E-6   -5.318909E-5   5.412092E-5   -1.693525E+2   -7.935250E+1   
5.073630E+3   1.399955E+2   1.399955E+2   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   -3.216033E-2   4.996979E-2   -5.242782E-5   -8.882059E-6   8.882059E-6   -5.242782E-5   5.317487E-5   -1.703845E+2   -8.038453E+1   
5.095909E+3   1.401039E+2   1.401039E+2   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   -3.102763E-2   5.283770E-2   -5.359537E-5   -1.159480E-5   1.159480E-5   -5.359537E-5   5.483523E-5   -1.677928E+2   -7.779278E+1   
5.118148E+3   1.399733E+2   1.399733E+2   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   -3.110985E-2   5.187990E-2   -5.302239E-5   -1.090780E-5   1.090780E-5   -5.302239E-5   5.413275E-5   -1.683753E+2   -7.837525E+1   
5.140462E+3   1.400239E+2   1.400239E+2   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   -3.174156E-2   5.102884E-2   -5.285866E-5   -9.884171E-6   9.884171E-6   -5.285866E-5   5.377485E-5   -1.694084E+2   -7.940844E+1   
5.162698E+3   1.401027E+2   1.401027E+2   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   -3.107395E-2   5.167588E-2   -5.286732E-5   -1.080097E-5   1.080097E-5   -5.286732E-5   5.395938E-5   -1.684532E+2   -7.845319E+1   
5.184916E+3   1.400112E+2   1.400112E+2   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   -3.134549E-2   5.156881E-2   -5.296546E-5   -1.053013E-5   1.053013E-5   -5.296546E-5   5.400207E-5   -1.687556E+2   -7.875557E+1   
5.207154E+3   1.400122E+2   1.400122E+2   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   -3.231585E-2   5.197868E-2   -5.383234E-5   -1.008039E-5   1.008039E-5   -5.383234E-5   5.476801E-5   -1.693939E+2   -7.939389E+1   
5.229341E+3   1.399957E+2   1.399957E+2   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   -3.132215E-2   5.176086E-2   -5.307612E-5   -1.067295E-5   1.067295E-5   -5.307612E-5   5.413858E-5   -1.686302E+2   -7.863016E+1   
5.251630E+3   1.400576E+2   1.400576E+2   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   -3.386762E-2   5.156144E-2   -5.451997E-5   -8.659871E-6   8.659871E-6   -5.451997E-5   5.520345E-5   -1.709746E+2   -8.097462E+1   
5.273902E+3   1.401251E+2   1.401251E+2   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   -3.237568E-2   5.157280E-2   -5.360498E-5   -9.770781E-6   9.770781E-6   -5.360498E-5   5.448818E-5   -1.696699E+2   -7.966989E+1   
5.296137E+3   1.400646E+2   1.400646E+2   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   -3.243000E-2   5.092393E-2   -5.321596E-5   -9.306388E-6   9.306388E-6   -5.321596E-5   5.402358E-5   -1.700804E+2   -8.008044E+1   
5.318409E+3   1.399928E+2   1.399928E+2   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   -3.268095E-2   5.119298E-2   -5.354634E-5   -9.296676E-6   9.296676E-6   -5.354634E-5   5.434739E-5   -1.701505E+2   -8.015053E+1   
5.340690E+3   1.400283E+2   1.400283E+2   -1.500000E+1   -1.500000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   -3.278250E-2   5.148443E-2   -5.379894E-5   -9.412107E-6   9.412107E-6   -5.379894E-5   5.461605E-5   -1.700766E+2   -8.007655E+1   
5.361888E+3   1.400669E+2   1.400669E+2   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   -3.204526E-2   5.197225E-2   -5.366085E-5   -1.027632E-5   1.027632E-5   -5.366085E-5   5.463598E-5   -1.691588E+2   -7.915883E+1   
5.384083E+3   1.400403E+2   1.400403E+2   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   -3.225176E-2   5.181545E-2   -5.368640E-5   -1.002108E-5   1.002108E-5   -5.368640E-5   5.461366E-5   -1.694269E+2   -7.942687E+1   
5.406267E+3   1.401006E+2   1.401006E+2   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   -3.288835E-2   5.171914E-2   -5.401724E-5   -9.487270E-6   9.487270E-6   -5.401724E-5   5.484406E-5   -1.700385E+2   -8.003851E+1   
5.428346E+3   1.399846E+2   1.399846E+2   -7.000000E+0   -7.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   -3.199128E-2   5.264872E-2   -5.406806E-5   -1.075850E-5   1.075850E-5   -5.406806E-5   5.512803E-5   -1.687462E+2   -7.874623E+1   
5.449438E+3   1.400143E+2   1.400143E+2   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   -3.190016E-2   5.241308E-2   -5.385826E-5   -1.067184E-5   1.067184E-5   -5.385826E-5   5.490538E-5   -1.687922E+2   -7.879220E+1   
5.471546E+3   1.400296E+2   1.400296E+2   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   -3.278925E-2   5.280274E-2   -5.466171E-5   -1.026899E-5   1.026899E-5   -5.466171E-5   5.561793E-5   -1.693602E+2   -7.936017E+1   
5.493663E+3   1.400428E+2   1.400428E+2   -1.000000E+0   -1.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   -3.303223E-2   5.286684E-2   -5.485369E-5   -1.013118E-5   1.013118E-5   -5.485369E-5   5.578143E-5   -1.695357E+2   -7.953570E+1   
5.514696E+3   1.400503E+2   1.400503E+2   0.000000E+0   0.000000E+0   9.000000E+1   0.000000E+0   0.000000E+0   -3.394218E-2   5.245698E-2   -5.514932E-5   -9.190201E-6   9.190201E-6   -5.514932E-5   5.590982E-5   -1.705390E+2   -8.053905E+1   
5.536647E+3   1.401211E+2   1.401211E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   -3.348014E-2   5.298559E-2   -5.520794E-5   -9.877531E-6   9.877531E-6   -5.520794E-5   5.608459E-5   -1.698562E+2   -7.985625E+1   
5.558158E+3   1.400541E+2   1.400541E+2   3.000000E+0   3.000000E+0   9.000000E+1   4.000000E+0   4.000000E+0   -3.305031E-2   5.134420E-2   -5.387319E-5   -9.122351E-6   9.122351E-6   -5.387319E-5   5.464007E-5   -1.703893E+2   -8.038926E+1   
5.579841E+3   1.399859E+2   1.399859E+2   5.000000E+0   5.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   -3.308777E-2   5.278033E-2   -5.483168E-5   -1.003355E-5   1.003355E-5   -5.483168E-5   5.574213E-5   -1.696303E+2   -7.963028E+1   
5.601489E+3   1.400456E+2   1.400456E+2   7.000000E+0   7.000000E+0   9.000000E+1   8.000000E+0   8.000000E+0   -3.227292E-2   5.302423E-2   -5.448675E-5   -1.079569E-5   1.079569E-5   -5.448675E-5   5.554595E-5   -1.687929E+2   -7.879290E+1   
5.623240E+3   1.400588E+2   1.400588E+2   9.000000E+0   9.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   -3.211767E-2   5.249502E-2   -5.404609E-5   -1.056454E-5   1.056454E-5   -5.404609E-5   5.506895E-5   -1.689397E+2   -7.893970E+1   
5.645274E+3   1.400193E+2   1.400193E+2   1.100000E+1   1.100000E+1   9.000000E+1   1.100000E+1   1.100000E+1   -3.205448E-2   5.301750E-2   -5.434731E-5   -1.095285E-5   1.095285E-5   -5.434731E-5   5.544001E-5   -1.686056E+2   -7.860556E+1   
5.667321E+3   1.400241E+2   1.400241E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   -3.374581E-2   5.276532E-2   -5.522873E-5   -9.537025E-6   9.537025E-6   -5.522873E-5   5.604612E-5   -1.702027E+2   -8.020265E+1   
5.689228E+3   1.400634E+2   1.400634E+2   1.500000E+1   1.500000E+1   9.000000E+1   1.500000E+1   1.500000E+1   -3.323869E-2   5.350959E-2   -5.539994E-5   -1.039869E-5   1.039869E-5   -5.539994E-5   5.636743E-5   -1.693692E+2   -7.936915E+1   
5.711308E+3   1.399915E+2   1.399915E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   -3.344518E-2   5.228792E-2   -5.473194E-5   -9.447274E-6   9.447274E-6   -5.473194E-5   5.554130E-5   -1.702067E+2   -8.020668E+1   
5.733162E+3   1.400180E+2   1.400180E+2   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   -3.352862E-2   5.346849E-2   -5.555242E-5   -1.015738E-5   1.015738E-5   -5.555242E-5   5.647339E-5   -1.696383E+2   -7.963832E+1   
5.755043E+3   1.400120E+2   1.400120E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   -3.373141E-2   5.282606E-2   -5.525939E-5   -9.587384E-6   9.587384E-6   -5.525939E-5   5.608492E-5   -1.701573E+2   -8.015729E+1   
5.776889E+3   1.400388E+2   1.400388E+2   2.300000E+1   2.300000E+1   9.000000E+1   2.300000E+1   2.300000E+1   -3.220236E-2   5.428760E-2   -5.526594E-5   -1.167384E-5   1.167384E-5   -5.526594E-5   5.648542E-5   -1.680727E+2   -7.807273E+1   
5.798974E+3   1.399812E+2   1.399812E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   -3.451895E-2   5.237689E-2   -5.545374E-5   -8.711247E-6   8.711247E-6   -5.545374E-5   5.613380E-5   -1.710723E+2   -8.107235E+1   
5.820907E+3   1.400547E+2   1.400547E+2   2.700000E+1   2.700000E+1   9.000000E+1   2.800000E+1   2.800000E+1   -3.335221E-2   5.340313E-2   -5.540079E-5   -1.024513E-5   1.024513E-5   -5.540079E-5   5.634013E-5   -1.695228E+2   -7.952280E+1   
5.842979E+3   1.400601E+2   1.400601E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   -3.265548E-2   5.425018E-2   -5.552171E-5   -1.131423E-5   1.131423E-5   -5.552171E-5   5.666280E-5   -1.684820E+2   -7.848196E+1   
5.864915E+3   1.400246E+2   1.400246E+2   3.100000E+1   3.100000E+1   9.000000E+1   3.100000E+1   3.100000E+1   -3.408790E-2   5.348138E-2   -5.590659E-5   -9.752142E-6   9.752142E-6   -5.590659E-5   5.675078E-5   -1.701051E+2   -8.010509E+1   
5.886998E+3   1.400698E+2   1.400698E+2   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   -3.395353E-2   5.336755E-2   -5.574938E-5   -9.777109E-6   9.777109E-6   -5.574938E-5   5.660022E-5   -1.700528E+2   -8.005285E+1   
5.908892E+3   1.400118E+2   1.400118E+2   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   -3.414833E-2   5.330310E-2   -5.582783E-5   -9.590896E-6   9.590896E-6   -5.582783E-5   5.664567E-5   -1.702521E+2   -8.025207E+1   
5.930783E+3   1.400105E+2   1.400105E+2   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   -3.252909E-2   5.340804E-2   -5.489510E-5   -1.085714E-5   1.085714E-5   -5.489510E-5   5.595846E-5   -1.688124E+2   -7.881243E+1   
5.952718E+3   1.400421E+2   1.400421E+2   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   -3.369121E-2   5.242845E-2   -5.497558E-5   -9.357175E-6   9.357175E-6   -5.497558E-5   5.576622E-5   -1.703405E+2   -8.034048E+1   
5.974556E+3   1.400081E+2   1.400081E+2   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   -3.381209E-2   5.310400E-2   -5.549028E-5   -9.709423E-6   9.709423E-6   -5.549028E-5   5.633333E-5   -1.700751E+2   -8.007513E+1   
5.996444E+3   1.400340E+2   1.400340E+2   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   -3.312550E-2   5.356971E-2   -5.536911E-5   -1.052171E-5   1.052171E-5   -5.536911E-5   5.635996E-5   -1.692405E+2   -7.924045E+1   
6.018384E+3   1.401062E+2   1.401062E+2   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   -3.375596E-2   5.308222E-2   -5.544140E-5   -9.736705E-6   9.736705E-6   -5.544140E-5   5.628989E-5   -1.700392E+2   -8.003920E+1   
6.040312E+3   1.399262E+2   1.399262E+2   4.700000E+1   4.700000E+1   9.000000E+1   4.700000E+1   4.700000E+1   -3.403697E-2   5.314573E-2   -5.565650E-5   -9.570377E-6   9.570377E-6   -5.565650E-5   5.647334E-5   -1.702432E+2   -8.024316E+1   
6.062336E+3   1.399803E+2   1.399803E+2   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   -3.469198E-2   5.335618E-2   -5.619852E-5   -9.223500E-6   9.223500E-6   -5.619852E-5   5.695039E-5   -1.706795E+2   -8.067951E+1   
6.096228E+3   1.399730E+2   1.399730E+2   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   -3.451619E-2   5.556662E-2   -5.752947E-5   -1.079864E-5   1.079864E-5   -5.752947E-5   5.853418E-5   -1.693689E+2   -7.936893E+1   
6.118829E+3   1.400824E+2   1.400824E+2   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   -3.602561E-2   5.649990E-2   -5.907050E-5   -1.029238E-5   1.029238E-5   -5.907050E-5   5.996046E-5   -1.701161E+2   -8.011607E+1   
6.141193E+3   1.400471E+2   1.400471E+2   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   -3.677541E-2   5.848730E-2   -6.082843E-5   -1.103711E-5   1.103711E-5   -6.082843E-5   6.182165E-5   -1.697158E+2   -7.971577E+1   
6.163572E+3   1.400229E+2   1.400229E+2   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   -3.760743E-2   5.961046E-2   -6.207433E-5   -1.115601E-5   1.115601E-5   -6.207433E-5   6.306885E-5   -1.698116E+2   -7.981155E+1   
6.186157E+3   1.400511E+2   1.400511E+2   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   -3.790655E-2   6.203105E-2   -6.383577E-5   -1.251729E-5   1.251729E-5   -6.383577E-5   6.505142E-5   -1.689059E+2   -7.890587E+1   
6.208531E+3   1.400727E+2   1.400727E+2   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   -3.958533E-2   6.330238E-2   -6.570167E-5   -1.210677E-5   1.210677E-5   -6.570167E-5   6.680781E-5   -1.695593E+2   -7.955930E+1   
6.230922E+3   1.400136E+2   1.400136E+2   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   -4.056154E-2   6.470169E-2   -6.721657E-5   -1.229956E-5   1.229956E-5   -6.721657E-5   6.833261E-5   -1.696305E+2   -7.963050E+1   
6.253504E+3   1.400885E+2   1.400885E+2   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   -4.108737E-2   6.629147E-2   -6.857706E-5   -1.295000E-5   1.295000E-5   -6.857706E-5   6.978908E-5   -1.693063E+2   -7.930627E+1   
6.275906E+3   1.399784E+2   1.399784E+2   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   -4.222926E-2   6.662373E-2   -6.949943E-5   -1.232264E-5   1.232264E-5   -6.949943E-5   7.058341E-5   -1.699456E+2   -7.994563E+1   
6.298095E+3   1.400549E+2   1.400549E+2   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   -4.420778E-2   6.881760E-2   -7.215149E-5   -1.229356E-5   1.229356E-5   -7.215149E-5   7.319132E-5   -1.703305E+2   -8.033049E+1   
6.321387E+3   1.400410E+2   1.400410E+2   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   -4.521500E-2   7.046539E-2   -7.384739E-5   -1.262586E-5   1.262586E-5   -7.384739E-5   7.491895E-5   -1.702978E+2   -8.029782E+1   
6.344004E+3   1.399907E+2   1.399907E+2   6.480000E+2   6.480000E+2   9.000000E+1   6.480000E+2   6.480000E+2   -4.678457E-2   7.229448E-2   -7.600904E-5   -1.266076E-5   1.266076E-5   -7.600904E-5   7.705627E-5   -1.705431E+2   -8.054311E+1   
6.366661E+3   1.400762E+2   1.400762E+2   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   -4.671710E-2   7.255004E-2   -7.613376E-5   -1.287775E-5   1.287775E-5   -7.613376E-5   7.721520E-5   -1.703995E+2   -8.039950E+1   
6.390041E+3   1.400810E+2   1.400810E+2   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   -4.813208E-2   7.530227E-2   -7.880107E-5   -1.363052E-5   1.363052E-5   -7.880107E-5   7.997124E-5   -1.701864E+2   -8.018644E+1   
6.412700E+3   1.400593E+2   1.400593E+2   7.980000E+2   7.980000E+2   9.000000E+1   7.980000E+2   7.980000E+2   -4.804126E-2   7.733446E-2   -8.006847E-5   -1.502628E-5   1.502628E-5   -8.006847E-5   8.146624E-5   -1.693710E+2   -7.937105E+1   
6.435303E+3   1.399945E+2   1.399945E+2   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   -4.863921E-2   7.844600E-2   -8.116208E-5   -1.531070E-5   1.531070E-5   -8.116208E-5   8.259359E-5   -1.693171E+2   -7.931706E+1   
6.458579E+3   1.401175E+2   1.401175E+2   8.980000E+2   8.980000E+2   9.000000E+1   8.980000E+2   8.980000E+2   -4.924390E-2   7.938047E-2   -8.214454E-5   -1.547440E-5   1.547440E-5   -8.214454E-5   8.358937E-5   -1.693316E+2   -7.933164E+1   
6.481211E+3   1.400639E+2   1.400639E+2   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   -5.098313E-2   8.079479E-2   -8.414094E-5   -1.511264E-5   1.511264E-5   -8.414094E-5   8.548737E-5   -1.698176E+2   -7.981761E+1   
6.503848E+3   1.400428E+2   1.400428E+2   9.980000E+2   9.980000E+2   9.000000E+1   9.980000E+2   9.980000E+2   -5.253092E-2   8.269414E-2   -8.633489E-5   -1.520959E-5   1.520959E-5   -8.633489E-5   8.766438E-5   -1.700087E+2   -8.000874E+1   
6.527324E+3   1.400665E+2   1.400665E+2   1.048000E+3   1.048000E+3   9.000000E+1   1.048000E+3   1.048000E+3   -5.447566E-2   8.378172E-2   -8.824555E-5   -1.448223E-5   1.448223E-5   -8.824555E-5   8.942601E-5   -1.706801E+2   -8.068010E+1   
6.550084E+3   1.400098E+2   1.400098E+2   1.098000E+3   1.098000E+3   9.000000E+1   1.098000E+3   1.098000E+3   -5.389154E-2   8.547858E-2   -8.898956E-5   -1.602363E-5   1.602363E-5   -8.898956E-5   9.042068E-5   -1.697926E+2   -7.979259E+1   
6.572882E+3   1.400082E+2   1.400082E+2   1.147000E+3   1.147000E+3   9.000000E+1   1.148000E+3   1.148000E+3   -5.491562E-2   8.731322E-2   -9.081758E-5   -1.646562E-5   1.646562E-5   -9.081758E-5   9.229815E-5   -1.697237E+2   -7.972366E+1   
6.596173E+3   1.400693E+2   1.400693E+2   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   -5.533561E-2   8.913680E-2   -9.226491E-5   -1.734719E-5   1.734719E-5   -9.226491E-5   9.388152E-5   -1.693518E+2   -7.935184E+1   
6.619008E+3   1.400900E+2   1.400900E+2   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   -5.619585E-2   8.996975E-2   -9.333925E-5   -1.725548E-5   1.725548E-5   -9.333925E-5   9.492085E-5   -1.695261E+2   -7.952607E+1   
6.642062E+3   1.399845E+2   1.399845E+2   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   -5.891035E-2   9.194739E-2   -9.630549E-5   -1.654068E-5   1.654068E-5   -9.630549E-5   9.771562E-5   -1.702544E+2   -8.025441E+1   
6.665306E+3   1.400730E+2   1.400730E+2   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   -5.938896E-2   9.343941E-2   -9.757313E-5   -1.716213E-5   1.716213E-5   -9.757313E-5   9.907096E-5   -1.700243E+2   -8.002429E+1   
6.687888E+3   1.400586E+2   1.400586E+2   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   -6.053207E-2   9.434569E-2   -9.887010E-5   -1.690915E-5   1.690915E-5   -9.887010E-5   1.003056E-4   -1.702949E+2   -8.029495E+1   
6.710427E+3   1.399855E+2   1.399855E+2   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   -6.160645E-2   9.751442E-2   -1.015981E-4   -1.818613E-5   1.818613E-5   -1.015981E-4   1.032129E-4   -1.698515E+2   -7.985149E+1   
6.733234E+3   1.399607E+2   1.399607E+2   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   -6.146349E-2   9.896676E-2   -1.024556E-4   -1.924136E-5   1.924136E-5   -1.024556E-4   1.042467E-4   -1.693636E+2   -7.936363E+1   
6.755751E+3   1.400735E+2   1.400735E+2   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   -6.282411E-2   9.900542E-2   -1.033220E-4   -1.826028E-5   1.826028E-5   -1.033220E-4   1.049232E-4   -1.699775E+2   -7.997751E+1   
6.778385E+3   1.400256E+2   1.400256E+2   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   -6.322724E-2   1.014217E-1   -1.051449E-4   -1.954183E-5   1.954183E-5   -1.051449E-4   1.069455E-4   -1.694714E+2   -7.947136E+1   
6.801415E+3   1.399848E+2   1.399848E+2   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   -6.505543E-2   1.021000E-1   -1.067170E-4   -1.863311E-5   1.863311E-5   -1.067170E-4   1.083315E-4   -1.700958E+2   -8.009583E+1   
6.823941E+3   1.400673E+2   1.400673E+2   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   -6.498701E-2   1.034561E-1   -1.075579E-4   -1.957024E-5   1.957024E-5   -1.075579E-4   1.093238E-4   -1.696878E+2   -7.968780E+1   
6.846504E+3   1.399780E+2   1.399780E+2   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   -6.702073E-2   1.053020E-1   -1.100175E-4   -1.927289E-5   1.927289E-5   -1.100175E-4   1.116928E-4   -1.700637E+2   -8.006373E+1   
6.869280E+3   1.400027E+2   1.400027E+2   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   -6.628841E-2   1.068716E-1   -1.105869E-4   -2.084067E-5   2.084067E-5   -1.105869E-4   1.125336E-4   -1.693275E+2   -7.932749E+1   
6.891819E+3   1.400427E+2   1.400427E+2   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   -6.964075E-2   1.087495E-1   -1.138826E-4   -1.958888E-5   1.958888E-5   -1.138826E-4   1.155550E-4   -1.702401E+2   -8.024009E+1   
6.914317E+3   1.399672E+2   1.399672E+2   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   -7.038592E-2   1.111320E-1   -1.158950E-4   -2.059536E-5   2.059536E-5   -1.158950E-4   1.177107E-4   -1.699233E+2   -7.992333E+1   
6.937088E+3   1.401089E+2   1.401089E+2   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   -7.006964E-2   1.120923E-1   -1.163248E-4   -2.145708E-5   2.145708E-5   -1.163248E-4   1.182872E-4   -1.695488E+2   -7.954880E+1   
6.959669E+3   1.399781E+2   1.399781E+2   1.999000E+3   1.999000E+3   9.000000E+1   2.000000E+3   2.000000E+3   -7.184781E-2   1.139705E-1   -1.186474E-4   -2.136980E-5   2.136980E-5   -1.186474E-4   1.205565E-4   -1.697898E+2   -7.978982E+1   
6.997561E+3   1.399894E+2   1.399894E+2   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   -8.121510E-2   1.289852E-1   -1.342177E-4   -2.425767E-5   2.425767E-5   -1.342177E-4   1.363921E-4   -1.697553E+2   -7.975531E+1   
7.024454E+3   1.400884E+2   1.400884E+2   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   -9.161145E-2   1.435876E-1   -1.501556E-4   -2.611485E-5   2.611485E-5   -1.501556E-4   1.524096E-4   -1.701339E+2   -8.013388E+1   
7.050405E+3   1.400680E+2   1.400680E+2   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -1.002081E-1   1.596909E-1   -1.659583E-4   -3.028438E-5   3.028438E-5   -1.659583E-4   1.686988E-4   -1.696583E+2   -7.965835E+1   
7.076259E+3   1.400558E+2   1.400558E+2   3.999000E+3   3.999000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -1.055696E-1   1.680476E-1   -1.747157E-4   -3.178221E-5   3.178221E-5   -1.747157E-4   1.775829E-4   -1.696902E+2   -7.969016E+1   
7.102612E+3   1.399842E+2   1.399842E+2   4.498000E+3   4.498000E+3   9.000000E+1   4.499000E+3   4.499000E+3   -1.036159E-1   1.686148E-1   -1.738772E-4   -3.359806E-5   3.359806E-5   -1.738772E-4   1.770936E-4   -1.690636E+2   -7.906360E+1   
7.128521E+3   1.400308E+2   1.400308E+2   4.997000E+3   4.997000E+3   9.000000E+1   4.999000E+3   4.999000E+3   -8.760166E-2   1.574399E-1   -1.566984E-4   -3.813687E-5   3.813687E-5   -1.566984E-4   1.612725E-4   -1.663214E+2   -7.632143E+1   
7.154200E+3   1.399371E+2   1.399371E+2   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -7.020096E-2   1.387826E-1   -1.337892E-4   -3.880935E-5   3.880935E-5   -1.337892E-4   1.393044E-4   -1.638237E+2   -7.382370E+1   
7.180621E+3   1.400250E+2   1.400250E+2   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -5.290673E-2   1.214482E-1   -1.118074E-4   -4.026796E-5   4.026796E-5   -1.118074E-4   1.188377E-4   -1.601933E+2   -7.019327E+1   
7.206607E+3   1.399878E+2   1.399878E+2   6.498000E+3   6.498000E+3   9.000000E+1   6.499000E+3   6.499000E+3   -4.547856E-2   1.164659E-1   -1.039700E-4   -4.250478E-5   4.250478E-5   -1.039700E-4   1.123228E-4   -1.577644E+2   -6.776439E+1   
7.232800E+3   1.399874E+2   1.399874E+2   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -4.547765E-2   1.197173E-1   -1.060870E-4   -4.463111E-5   4.463111E-5   -1.060870E-4   1.150930E-4   -1.571834E+2   -6.718337E+1   
7.258464E+3   1.400341E+2   1.400341E+2   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -4.972126E-2   1.292687E-1   -1.149313E-4   -4.773683E-5   4.773683E-5   -1.149313E-4   1.244509E-4   -1.574444E+2   -6.744440E+1   
7.283711E+3   1.400114E+2   1.400114E+2   7.999000E+3   7.999000E+3   9.000000E+1   8.000000E+3   8.000000E+3   -5.681251E-2   1.400126E-1   -1.263129E-4   -4.951597E-5   4.951597E-5   -1.263129E-4   1.356715E-4   -1.585943E+2   -6.859430E+1   
7.310121E+3   1.400744E+2   1.400744E+2   8.498000E+3   8.498000E+3   9.000000E+1   8.499000E+3   8.499000E+3   -6.402643E-2   1.523772E-1   -1.388258E-4   -5.226399E-5   5.226399E-5   -1.388258E-4   1.483379E-4   -1.593701E+2   -6.937006E+1   
7.336523E+3   1.399987E+2   1.399987E+2   8.998000E+3   8.998000E+3   9.000000E+1   8.999000E+3   8.999000E+3   -7.336153E-2   1.676785E-1   -1.545628E-4   -5.536300E-5   5.536300E-5   -1.545628E-4   1.641789E-4   -1.602929E+2   -7.029293E+1   
7.362951E+3   1.399978E+2   1.399978E+2   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -8.705524E-2   1.869941E-1   -1.756089E-4   -5.786271E-5   5.786271E-5   -1.756089E-4   1.848961E-4   -1.617631E+2   -7.176307E+1   
7.388211E+3   1.400105E+2   1.400105E+2   9.998000E+3   9.998000E+3   9.000000E+1   1.000000E+4   1.000000E+4   -1.023298E-1   2.080237E-1   -1.987487E-4   -6.031370E-5   6.031370E-5   -1.987487E-4   2.076988E-4   -1.631187E+2   -7.311868E+1   
@@END Data.
@Time at end of measurement: 12:49:45
@Instrument  Changes:
@Emu Range: 20 uV
@END Instrument  Changes:
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -9499.000      -9999.000      250.000        Coercive Field: Field at which M//H changes sign
Ms  emu                                 3.017E-4       -1.987E-4      2.502E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -5.515E-5      1.647E-4       1.099E-4       Remanent Magnetization: M at H=0        
S                                       0.183          0.829          0.506          Squareness: Mr/Ms                       
S*                                      1.372          1.151          1.261          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
