@Filename: c:\vsm-lv\Will\data\AJA335e-FePtFeRh_1030nm_Tann_6\AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_160deg.VHD
@Measurement Controlfilename: C:\vsm-lv\Will\Recipes\10kOe OoP loop 160deg.VHC
@Signal Manipulation filename: c:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA335e-FePtFeRh_1030nm_Tann_6
@Date: 12 November 2019    (2019-12-11)
@Time: 15:11:29
@Test ID: AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_160deg
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 90.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Sample Temperature to 160.0558 [degC] and wait 60.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Applied Field to 9999.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 3:      Set Auto Range Signal to 11.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 5
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 5.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 10000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To: 50.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: 50.0000 [Oe] To: -50.0000 [Oe] Min Stepsize/Sweeprate =  2.0000 [Oe] Max Stepsize/Sweeprate =  2.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -50.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -10000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 4 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 10 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.706
@Y Coils Correction Factor: 0.964
@Sample Shape Correction Factor: 0.919
@Coil Angle Alpha: 42.300
@Coil Angle Beta: -47.320
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
15000.000000   1.000000
15249.000000   1.000524
15499.000000   1.000702
15750.000000   1.001233
16000.000000   1.001406
16250.000000   1.001585
16499.000000   1.001758
16749.000000   1.001937
16999.000000   1.002110
17249.000000   1.001937
17499.000000   1.002289
17749.000000   1.002289
17999.000000   1.002289
18249.000000   1.002462
18499.000000   1.002462
18748.000000   1.002462
18999.000000   1.002462
19249.000000   1.002462
19499.000000   1.002642
19749.000000   1.002642
19999.000000   1.002462
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = No
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 25 October 2019  12:02:56
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 5
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 15:11:29
@@Data
New Section: Section 0: 
2.965900E+1   1.599936E+2   1.599936E+2   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -8.249811E-2   1.999320E-1   -1.812178E-4   -6.969173E-5   6.969173E-5   -1.812178E-4   1.941567E-4   -1.589645E+2   -6.896453E+1   
5.495700E+1   1.601221E+2   1.601221E+2   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -6.913884E-2   1.791452E-1   -1.594202E-4   -6.598281E-5   6.598281E-5   -1.594202E-4   1.725356E-4   -1.575157E+2   -6.751571E+1   
8.009800E+1   1.600542E+2   1.600542E+2   8.998000E+3   8.998000E+3   9.000000E+1   8.998000E+3   8.998000E+3   -5.978134E-2   1.643377E-1   -1.439910E-4   -6.322319E-5   6.322319E-5   -1.439910E-4   1.572596E-4   -1.562948E+2   -6.629481E+1   
1.049970E+2   1.600954E+2   1.600954E+2   8.498000E+3   8.498000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -4.763843E-2   1.452685E-1   -1.240642E-4   -5.973761E-5   5.973761E-5   -1.240642E-4   1.376971E-4   -1.542889E+2   -6.428892E+1   
1.303960E+2   1.599799E+2   1.599799E+2   7.999000E+3   7.999000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -4.416041E-2   1.328778E-1   -1.138439E-4   -5.420934E-5   5.420934E-5   -1.138439E-4   1.260916E-4   -1.545375E+2   -6.453750E+1   
1.559430E+2   1.599626E+2   1.599626E+2   7.498000E+3   7.498000E+3   9.000000E+1   7.498000E+3   7.498000E+3   -2.855104E-2   1.112732E-1   -9.012261E-5   -5.163002E-5   5.163002E-5   -9.012261E-5   1.038641E-4   -1.501922E+2   -6.019219E+1   
1.812810E+2   1.600588E+2   1.600588E+2   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -1.764634E-2   9.490916E-2   -7.272312E-5   -4.899714E-5   4.899714E-5   -7.272312E-5   8.768907E-5   -1.460299E+2   -5.602991E+1   
2.066760E+2   1.600207E+2   1.600207E+2   6.498000E+3   6.498000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -9.042148E-3   7.746257E-2   -5.604083E-5   -4.395499E-5   4.395499E-5   -5.604083E-5   7.122230E-5   -1.418915E+2   -5.189154E+1   
2.319850E+2   1.601081E+2   1.601081E+2   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -3.121325E-3   6.435270E-2   -4.384198E-5   -3.976335E-5   3.976335E-5   -4.384198E-5   5.918820E-5   -1.377929E+2   -4.779292E+1   
2.578200E+2   1.599823E+2   1.599823E+2   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   1.063027E-2   4.733960E-2   -2.425965E-5   -3.881177E-5   3.881177E-5   -2.425965E-5   4.576991E-5   -1.220078E+2   -3.200781E+1   
2.834000E+2   1.599643E+2   1.599643E+2   4.997000E+3   4.997000E+3   9.000000E+1   4.998000E+3   4.998000E+3   2.149860E-2   2.900066E-2   -5.596385E-6   -3.486085E-5   3.486085E-5   -5.596385E-6   3.530720E-5   -9.912016E+1   -9.120161E+0   
3.090210E+2   1.600103E+2   1.600103E+2   4.498000E+3   4.498000E+3   9.000000E+1   4.498000E+3   4.498000E+3   3.185124E-2   1.338666E-2   1.097333E-5   -3.230999E-5   3.230999E-5   1.097333E-5   3.412256E-5   -7.124114E+1   1.875886E+1   
3.352400E+2   1.600520E+2   1.600520E+2   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   4.095654E-2   -4.291133E-3   2.811602E-5   -2.748731E-5   2.748731E-5   2.811602E-5   3.932001E-5   -4.435218E+1   4.564782E+1   
3.610690E+2   1.599991E+2   1.599991E+2   3.498000E+3   3.498000E+3   9.000000E+1   3.498000E+3   3.498000E+3   5.059609E-2   -2.096584E-2   4.493570E-5   -2.371556E-5   2.371556E-5   4.493570E-5   5.080989E-5   -2.782360E+1   6.217640E+1   
3.864330E+2   1.600336E+2   1.600336E+2   2.998000E+3   2.998000E+3   9.000000E+1   2.998000E+3   2.998000E+3   6.165263E-2   -3.623178E-2   6.171391E-5   -2.191289E-5   2.191289E-5   6.171391E-5   6.548879E-5   -1.954853E+1   7.045147E+1   
4.120410E+2   1.600250E+2   1.600250E+2   2.498000E+3   2.498000E+3   9.000000E+1   2.498000E+3   2.498000E+3   7.245970E-2   -5.522455E-2   8.076514E-5   -1.748920E-5   1.748920E-5   8.076514E-5   8.263704E-5   -1.221840E+1   7.778160E+1   
4.374410E+2   1.599764E+2   1.599764E+2   1.998000E+3   1.998000E+3   9.000000E+1   1.999000E+3   1.999000E+3   8.275825E-2   -7.150910E-2   9.773814E-5   -1.445994E-5   1.445994E-5   9.773814E-5   9.880200E-5   -8.415622E+0   8.158438E+1   
4.713040E+2   1.600588E+2   1.600588E+2   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   8.297194E-2   -7.192557E-2   9.814150E-5   -1.434572E-5   1.434572E-5   9.814150E-5   9.918444E-5   -8.316246E+0   8.168375E+1   
4.935900E+2   1.600527E+2   1.600527E+2   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   8.261868E-2   -7.277770E-2   9.847808E-5   -1.352734E-5   1.352734E-5   9.847808E-5   9.940282E-5   -7.821426E+0   8.217857E+1   
5.158470E+2   1.600144E+2   1.600144E+2   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   8.624359E-2   -7.475420E-2   1.020064E-4   -1.491625E-5   1.491625E-5   1.020064E-4   1.030913E-4   -8.319316E+0   8.168068E+1   
5.380950E+2   1.599973E+2   1.599973E+2   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   8.597943E-2   -7.757960E-2   1.036833E-4   -1.287371E-5   1.287371E-5   1.036833E-4   1.044794E-4   -7.077838E+0   8.292216E+1   
5.601400E+2   1.599924E+2   1.599924E+2   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   8.600858E-2   -7.942541E-2   1.049035E-4   -1.168853E-5   1.168853E-5   1.049035E-4   1.055526E-4   -6.357773E+0   8.364223E+1   
5.823960E+2   1.600306E+2   1.600306E+2   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   8.779459E-2   -8.061286E-2   1.067810E-4   -1.223319E-5   1.223319E-5   1.067810E-4   1.074795E-4   -6.535503E+0   8.346450E+1   
6.046810E+2   1.600106E+2   1.600106E+2   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   8.878261E-2   -8.026067E-2   1.071625E-4   -1.319422E-5   1.319422E-5   1.071625E-4   1.079717E-4   -7.019128E+0   8.298087E+1   
6.267190E+2   1.600164E+2   1.600164E+2   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   8.924787E-2   -8.268095E-2   1.090264E-4   -1.195603E-5   1.195603E-5   1.090264E-4   1.096800E-4   -6.258149E+0   8.374185E+1   
6.487540E+2   1.600386E+2   1.600386E+2   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   9.130233E-2   -8.499495E-2   1.118037E-4   -1.196274E-5   1.196274E-5   1.118037E-4   1.124418E-4   -6.107283E+0   8.389272E+1   
6.707410E+2   1.600404E+2   1.600404E+2   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   9.119053E-2   -8.628621E-2   1.125755E-4   -1.103586E-5   1.103586E-5   1.125755E-4   1.131152E-4   -5.598856E+0   8.440114E+1   
6.930850E+2   1.599991E+2   1.599991E+2   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   9.159887E-2   -8.824049E-2   1.141008E-4   -1.006023E-5   1.006023E-5   1.141008E-4   1.145434E-4   -5.038719E+0   8.496128E+1   
7.150660E+2   1.601009E+2   1.601009E+2   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   9.348005E-2   -9.000087E-2   1.164104E-4   -1.030072E-5   1.030072E-5   1.164104E-4   1.168652E-4   -5.056721E+0   8.494328E+1   
7.373220E+2   1.600293E+2   1.600293E+2   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   9.443330E-2   -9.035001E-2   1.172271E-4   -1.077752E-5   1.077752E-5   1.172271E-4   1.177215E-4   -5.252843E+0   8.474716E+1   
7.595490E+2   1.601189E+2   1.601189E+2   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   9.578371E-2   -9.210019E-2   1.192019E-4   -1.063210E-5   1.063210E-5   1.192019E-4   1.196751E-4   -5.096958E+0   8.490304E+1   
7.818630E+2   1.599118E+2   1.599118E+2   1.248000E+3   1.248000E+3   9.000000E+1   1.248000E+3   1.248000E+3   9.704345E-2   -9.525938E-2   1.220382E-4   -9.498460E-6   9.498460E-6   1.220382E-4   1.224073E-4   -4.450464E+0   8.554954E+1   
8.041660E+2   1.598885E+2   1.598885E+2   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   9.801875E-2   -9.501728E-2   1.224835E-4   -1.037810E-5   1.037810E-5   1.224835E-4   1.229224E-4   -4.843137E+0   8.515686E+1   
8.264440E+2   1.600200E+2   1.600200E+2   1.148000E+3   1.148000E+3   9.000000E+1   1.149000E+3   1.149000E+3   9.815866E-2   -9.735672E-2   1.240937E-4   -8.952117E-6   8.952117E-6   1.240937E-4   1.244162E-4   -4.126169E+0   8.587383E+1   
8.486480E+2   1.600410E+2   1.600410E+2   1.098000E+3   1.098000E+3   9.000000E+1   1.099000E+3   1.099000E+3   9.795554E-2   -9.896940E-2   1.250184E-4   -7.747560E-6   7.747560E-6   1.250184E-4   1.252582E-4   -3.546162E+0   8.645384E+1   
8.709520E+2   1.599948E+2   1.599948E+2   1.048000E+3   1.048000E+3   9.000000E+1   1.048000E+3   1.048000E+3   1.002775E-1   -9.973436E-2   1.269522E-4   -8.964879E-6   8.964879E-6   1.269522E-4   1.272683E-4   -4.039304E+0   8.596070E+1   
8.930720E+2   1.600364E+2   1.600364E+2   9.980000E+2   9.980000E+2   9.000000E+1   9.990000E+2   9.990000E+2   1.015546E-1   -1.012751E-1   1.287452E-4   -8.902130E-6   8.902130E-6   1.287452E-4   1.290526E-4   -3.955441E+0   8.604456E+1   
9.149990E+2   1.601427E+2   1.601427E+2   9.480000E+2   9.480000E+2   9.000000E+1   9.480000E+2   9.480000E+2   1.027121E-1   -1.033935E-1   1.308405E-4   -8.373299E-6   8.373299E-6   1.308405E-4   1.311082E-4   -3.661720E+0   8.633828E+1   
9.368420E+2   1.600115E+2   1.600115E+2   8.980000E+2   8.980000E+2   9.000000E+1   8.980000E+2   8.980000E+2   1.042964E-1   -1.047819E-1   1.327242E-4   -8.637421E-6   8.637421E-6   1.327242E-4   1.330050E-4   -3.723442E+0   8.627656E+1   
9.587240E+2   1.600459E+2   1.600459E+2   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   1.041545E-1   -1.077647E-1   1.345792E-4   -6.582394E-6   6.582394E-6   1.345792E-4   1.347401E-4   -2.800159E+0   8.719984E+1   
9.806030E+2   1.599696E+2   1.599696E+2   7.970000E+2   7.970000E+2   9.000000E+1   7.980000E+2   7.980000E+2   1.052781E-1   -1.074735E-1   1.350842E-4   -7.603810E-6   7.603810E-6   1.350842E-4   1.352981E-4   -3.221745E+0   8.677825E+1   
1.002496E+3   1.599657E+2   1.599657E+2   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   1.067796E-1   -1.092640E-1   1.371786E-4   -7.543790E-6   7.543790E-6   1.371786E-4   1.373859E-4   -3.147666E+0   8.685233E+1   
1.024330E+3   1.600636E+2   1.600636E+2   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   1.078951E-1   -1.111644E-1   1.391060E-4   -7.126396E-6   7.126396E-6   1.391060E-4   1.392884E-4   -2.932698E+0   8.706730E+1   
1.046264E+3   1.600930E+2   1.600930E+2   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   1.076602E-1   -1.118576E-1   1.394122E-4   -6.499502E-6   6.499502E-6   1.394122E-4   1.395637E-4   -2.669239E+0   8.733076E+1   
1.068145E+3   1.600693E+2   1.600693E+2   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   1.086811E-1   -1.139080E-1   1.413788E-4   -5.914033E-6   5.914033E-6   1.413788E-4   1.415025E-4   -2.395350E+0   8.760465E+1   
1.089987E+3   1.598747E+2   1.598747E+2   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   1.091698E-1   -1.153047E-1   1.425906E-4   -5.362389E-6   5.362389E-6   1.425906E-4   1.426914E-4   -2.153701E+0   8.784630E+1   
1.111828E+3   1.600411E+2   1.600411E+2   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   1.104140E-1   -1.163368E-1   1.440320E-4   -5.607916E-6   5.607916E-6   1.440320E-4   1.441411E-4   -2.229697E+0   8.777030E+1   
1.133708E+3   1.599880E+2   1.599880E+2   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   1.125178E-1   -1.170149E-1   1.457744E-4   -6.720609E-6   6.720609E-6   1.457744E-4   1.459292E-4   -2.639628E+0   8.736037E+1   
1.155582E+3   1.600941E+2   1.600941E+2   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   1.119759E-1   -1.199078E-1   1.473234E-4   -4.428482E-6   4.428482E-6   1.473234E-4   1.473899E-4   -1.721770E+0   8.827823E+1   
1.177433E+3   1.600309E+2   1.600309E+2   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   1.127194E-1   -1.209233E-1   1.484445E-4   -4.314487E-6   4.314487E-6   1.484445E-4   1.485071E-4   -1.664813E+0   8.833519E+1   
1.199264E+3   1.600298E+2   1.600298E+2   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   1.129749E-1   -1.244508E-1   1.508999E-4   -2.197352E-6   2.197352E-6   1.508999E-4   1.509159E-4   -8.342624E-1   8.916574E+1   
1.221144E+3   1.600880E+2   1.600880E+2   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   1.152584E-1   -1.239685E-1   1.519975E-4   -4.201578E-6   4.201578E-6   1.519975E-4   1.520556E-4   -1.583390E+0   8.841661E+1   
1.243021E+3   1.600016E+2   1.600016E+2   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   1.143537E-1   -1.266138E-1   1.531610E-4   -1.802957E-6   1.802957E-6   1.531610E-4   1.531716E-4   -6.744343E-1   8.932557E+1   
1.264858E+3   1.600510E+2   1.600510E+2   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   1.156698E-1   -1.277735E-1   1.547300E-4   -2.018242E-6   2.018242E-6   1.547300E-4   1.547432E-4   -7.473028E-1   8.925270E+1   
1.286702E+3   1.600422E+2   1.600422E+2   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   1.170318E-1   -1.289795E-1   1.563575E-4   -2.237207E-6   2.237207E-6   1.563575E-4   1.563735E-4   -8.197479E-1   8.918025E+1   
1.308431E+3   1.600070E+2   1.600070E+2   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   1.177793E-1   -1.306453E-1   1.579046E-4   -1.701053E-6   1.701053E-6   1.579046E-4   1.579137E-4   -6.172045E-1   8.938280E+1   
1.341622E+3   1.601345E+2   1.601345E+2   4.700000E+1   4.700000E+1   9.000000E+1   4.800000E+1   4.800000E+1   1.182860E-1   -1.306368E-1   1.582123E-4   -2.081306E-6   2.081306E-6   1.582123E-4   1.582260E-4   -7.536910E-1   8.924631E+1   
1.362994E+3   1.600803E+2   1.600803E+2   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   1.194141E-1   -1.307868E-1   1.590074E-4   -2.817602E-6   2.817602E-6   1.590074E-4   1.590324E-4   -1.015171E+0   8.898483E+1   
1.382001E+3   1.600824E+2   1.600824E+2   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   1.189856E-1   -1.308866E-1   1.588075E-4   -2.435522E-6   2.435522E-6   1.588075E-4   1.588262E-4   -8.786373E-1   8.912136E+1   
1.404441E+3   1.599833E+2   1.599833E+2   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   1.181792E-1   -1.300326E-1   1.577528E-4   -2.397384E-6   2.397384E-6   1.577528E-4   1.577710E-4   -8.706625E-1   8.912934E+1   
1.423597E+3   1.600166E+2   1.600166E+2   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   1.179319E-1   -1.300846E-1   1.576338E-4   -2.180487E-6   2.180487E-6   1.576338E-4   1.576488E-4   -7.924999E-1   8.920750E+1   
1.445953E+3   1.600128E+2   1.600128E+2   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   1.191764E-1   -1.294403E-1   1.579836E-4   -3.522165E-6   3.522165E-6   1.579836E-4   1.580228E-4   -1.277169E+0   8.872283E+1   
1.465018E+3   1.600312E+2   1.600312E+2   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   1.186118E-1   -1.307155E-1   1.584650E-4   -2.270854E-6   2.270854E-6   1.584650E-4   1.584813E-4   -8.210105E-1   8.917899E+1   
1.487424E+3   1.599872E+2   1.599872E+2   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   1.195544E-1   -1.310229E-1   1.592480E-4   -2.767054E-6   2.767054E-6   1.592480E-4   1.592720E-4   -9.954574E-1   8.900454E+1   
1.506534E+3   1.600330E+2   1.600330E+2   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   1.197793E-1   -1.312757E-1   1.595517E-4   -2.768113E-6   2.768113E-6   1.595517E-4   1.595757E-4   -9.939431E-1   8.900606E+1   
1.528963E+3   1.600469E+2   1.600469E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   1.181887E-1   -1.317862E-1   1.589008E-4   -1.257935E-6   1.257935E-6   1.589008E-4   1.589057E-4   -4.535716E-1   8.954643E+1   
1.548042E+3   1.601129E+2   1.601129E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   1.179289E-1   -1.305609E-1   1.579421E-4   -1.866830E-6   1.866830E-6   1.579421E-4   1.579531E-4   -6.771881E-1   8.932281E+1   
1.570389E+3   1.600019E+2   1.600019E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   1.175464E-1   -1.301300E-1   1.574250E-4   -1.865679E-6   1.865679E-6   1.574250E-4   1.574361E-4   -6.789935E-1   8.932101E+1   
1.589456E+3   1.600312E+2   1.600312E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   1.185062E-1   -1.309841E-1   1.585747E-4   -2.017184E-6   2.017184E-6   1.585747E-4   1.585875E-4   -7.288042E-1   8.927120E+1   
1.611891E+3   1.599646E+2   1.599646E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   1.193180E-1   -1.322093E-1   1.598745E-4   -1.816614E-6   1.816614E-6   1.598745E-4   1.598848E-4   -6.510095E-1   8.934899E+1   
1.630945E+3   1.600417E+2   1.600417E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   1.193709E-1   -1.308720E-1   1.590362E-4   -2.730039E-6   2.730039E-6   1.590362E-4   1.590597E-4   -9.834510E-1   8.901655E+1   
1.653331E+3   1.599633E+2   1.599633E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   1.181952E-1   -1.315365E-1   1.587421E-4   -1.425984E-6   1.425984E-6   1.587421E-4   1.587485E-4   -5.146755E-1   8.948532E+1   
1.672359E+3   1.599776E+2   1.599776E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   1.211589E-1   -1.313342E-1   1.604427E-4   -3.750351E-6   3.750351E-6   1.604427E-4   1.604865E-4   -1.339046E+0   8.866095E+1   
1.694792E+3   1.599532E+2   1.599532E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   1.194199E-1   -1.315570E-1   1.595127E-4   -2.318373E-6   2.318373E-6   1.595127E-4   1.595295E-4   -8.326841E-1   8.916732E+1   
1.713863E+3   1.600807E+2   1.600807E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   1.189102E-1   -1.310677E-1   1.588788E-4   -2.261284E-6   2.261284E-6   1.588788E-4   1.588949E-4   -8.154221E-1   8.918458E+1   
1.736040E+3   1.600666E+2   1.600666E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   1.178785E-1   -1.323105E-1   1.590505E-4   -6.857470E-7   6.857470E-7   1.590505E-4   1.590520E-4   -2.470295E-1   8.975297E+1   
1.754765E+3   1.600385E+2   1.600385E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   1.192209E-1   -1.320820E-1   1.597315E-4   -1.828021E-6   1.828021E-6   1.597315E-4   1.597420E-4   -6.556836E-1   8.934432E+1   
1.776756E+3   1.600402E+2   1.600402E+2   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   1.189790E-1   -1.319488E-1   1.594953E-4   -1.736161E-6   1.736161E-6   1.594953E-4   1.595047E-4   -6.236598E-1   8.937634E+1   
1.795508E+3   1.600897E+2   1.600897E+2   5.000000E+0   5.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   1.183840E-1   -1.322349E-1   1.593137E-4   -1.109038E-6   1.109038E-6   1.593137E-4   1.593176E-4   -3.988494E-1   8.960115E+1   
1.817171E+3   1.600371E+2   1.600371E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   1.176814E-1   -1.322160E-1   1.588671E-4   -6.017313E-7   6.017313E-7   1.588671E-4   1.588682E-4   -2.170147E-1   8.978299E+1   
1.835943E+3   1.600660E+2   1.600660E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   1.200355E-1   -1.311320E-1   1.596164E-4   -3.051558E-6   3.051558E-6   1.596164E-4   1.596456E-4   -1.095251E+0   8.890475E+1   
1.858037E+3   1.600280E+2   1.600280E+2   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   1.198250E-1   -1.324558E-1   1.603485E-4   -2.030422E-6   2.030422E-6   1.603485E-4   1.603613E-4   -7.254725E-1   8.927453E+1   
1.880116E+3   1.600828E+2   1.600828E+2   -3.000000E+0   -3.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   1.202634E-1   -1.321835E-1   1.604422E-4   -2.532696E-6   2.532696E-6   1.604422E-4   1.604622E-4   -9.043803E-1   8.909562E+1   
1.901801E+3   1.600866E+2   1.600866E+2   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   1.179623E-1   -1.312294E-1   1.583981E-4   -1.454509E-6   1.454509E-6   1.583981E-4   1.584048E-4   -5.261104E-1   8.947389E+1   
1.923873E+3   1.600109E+2   1.600109E+2   -7.000000E+0   -7.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   1.188466E-1   -1.332249E-1   1.602445E-4   -8.039713E-7   8.039713E-7   1.602445E-4   1.602466E-4   -2.874593E-1   8.971254E+1   
1.945594E+3   1.600858E+2   1.600858E+2   -9.000000E+0   -9.000000E+0   9.000000E+1   -9.000000E+0   -9.000000E+0   1.194125E-1   -1.331192E-1   1.605256E-4   -1.291611E-6   1.291611E-6   1.605256E-4   1.605308E-4   -4.609998E-1   8.953900E+1   
1.967424E+3   1.600285E+2   1.600285E+2   -1.100000E+1   -1.100000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   1.194375E-1   -1.321722E-1   1.599242E-4   -1.929278E-6   1.929278E-6   1.599242E-4   1.599358E-4   -6.911659E-1   8.930883E+1   
1.989312E+3   1.600387E+2   1.600387E+2   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   1.185059E-1   -1.322558E-1   1.594027E-4   -1.185582E-6   1.185582E-6   1.594027E-4   1.594071E-4   -4.261383E-1   8.957386E+1   
2.011531E+3   1.600933E+2   1.600933E+2   -1.500000E+1   -1.500000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   1.197708E-1   -1.327347E-1   1.604966E-4   -1.808054E-6   1.808054E-6   1.604966E-4   1.605068E-4   -6.454309E-1   8.935457E+1   
2.033454E+3   1.599771E+2   1.599771E+2   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   1.198387E-1   -1.320508E-1   1.600932E-4   -2.305285E-6   2.305285E-6   1.600932E-4   1.601098E-4   -8.249818E-1   8.917502E+1   
2.055658E+3   1.600425E+2   1.600425E+2   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   1.196461E-1   -1.325437E-1   1.602951E-4   -1.840676E-6   1.840676E-6   1.602951E-4   1.603057E-4   -6.579009E-1   8.934210E+1   
2.077920E+3   1.601211E+2   1.601211E+2   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   1.185668E-1   -1.326480E-1   1.596958E-4   -9.741893E-7   9.741893E-7   1.596958E-4   1.596988E-4   -3.495160E-1   8.965048E+1   
2.100145E+3   1.600410E+2   1.600410E+2   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   1.184198E-1   -1.327138E-1   1.596477E-4   -8.223933E-7   8.223933E-7   1.596477E-4   1.596498E-4   -2.951451E-1   8.970485E+1   
2.122413E+3   1.599663E+2   1.599663E+2   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   1.195328E-1   -1.326614E-1   1.603017E-4   -1.679906E-6   1.679906E-6   1.603017E-4   1.603105E-4   -6.004179E-1   8.939958E+1   
2.144676E+3   1.599896E+2   1.599896E+2   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   1.193104E-1   -1.328350E-1   1.602773E-4   -1.401875E-6   1.401875E-6   1.602773E-4   1.602834E-4   -5.011282E-1   8.949887E+1   
2.166950E+3   1.600966E+2   1.600966E+2   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   1.199491E-1   -1.318605E-1   1.600375E-4   -2.511412E-6   2.511412E-6   1.600375E-4   1.600572E-4   -8.990487E-1   8.910095E+1   
2.189188E+3   1.600688E+2   1.600688E+2   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   1.191915E-1   -1.329876E-1   1.603032E-4   -1.214167E-6   1.214167E-6   1.603032E-4   1.603078E-4   -4.339609E-1   8.956604E+1   
2.211412E+3   1.599810E+2   1.599810E+2   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   1.194274E-1   -1.330413E-1   1.604840E-4   -1.353556E-6   1.353556E-6   1.604840E-4   1.604897E-4   -4.832333E-1   8.951677E+1   
2.233604E+3   1.600302E+2   1.600302E+2   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   1.198212E-1   -1.333957E-1   1.609582E-4   -1.413153E-6   1.413153E-6   1.609582E-4   1.609644E-4   -5.030226E-1   8.949698E+1   
2.255872E+3   1.600595E+2   1.600595E+2   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   1.206840E-1   -1.339108E-1   1.618272E-4   -1.714587E-6   1.714587E-6   1.618272E-4   1.618362E-4   -6.070359E-1   8.939296E+1   
2.278159E+3   1.600630E+2   1.600630E+2   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   1.207233E-1   -1.330511E-1   1.612916E-4   -2.305606E-6   2.305606E-6   1.612916E-4   1.613080E-4   -8.189672E-1   8.918103E+1   
2.300399E+3   1.601119E+2   1.601119E+2   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   1.204900E-1   -1.328689E-1   1.610286E-4   -2.252198E-6   2.252198E-6   1.610286E-4   1.610444E-4   -8.013050E-1   8.919870E+1   
2.322680E+3   1.600853E+2   1.600853E+2   -4.300000E+1   -4.300000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   1.199110E-1   -1.333961E-1   1.610141E-4   -1.479332E-6   1.479332E-6   1.610141E-4   1.610209E-4   -5.263954E-1   8.947360E+1   
2.344571E+3   1.600532E+2   1.600532E+2   -4.500000E+1   -4.500000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   1.204777E-1   -1.323388E-1   1.606758E-4   -2.589703E-6   2.589703E-6   1.606758E-4   1.606966E-4   -9.233888E-1   8.907661E+1   
2.366501E+3   1.600657E+2   1.600657E+2   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.600000E+1   -4.600000E+1   1.202358E-1   -1.339956E-1   1.616053E-4   -1.327588E-6   1.327588E-6   1.616053E-4   1.616107E-4   -4.706743E-1   8.952933E+1   
2.388740E+3   1.600373E+2   1.600373E+2   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.800000E+1   -4.800000E+1   1.203596E-1   -1.343094E-1   1.618862E-4   -1.213976E-6   1.213976E-6   1.618862E-4   1.618908E-4   -4.296500E-1   8.957035E+1   
2.422059E+3   1.600193E+2   1.600193E+2   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   1.216687E-1   -1.346076E-1   1.628898E-4   -1.987253E-6   1.987253E-6   1.628898E-4   1.629019E-4   -6.989729E-1   8.930103E+1   
2.444488E+3   1.600505E+2   1.600505E+2   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   1.224780E-1   -1.365317E-1   1.646433E-4   -1.327954E-6   1.327954E-6   1.646433E-4   1.646486E-4   -4.621174E-1   8.953788E+1   
2.466129E+3   1.600514E+2   1.600514E+2   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   1.238546E-1   -1.373407E-1   1.660212E-4   -1.817213E-6   1.817213E-6   1.660212E-4   1.660312E-4   -6.271153E-1   8.937288E+1   
2.487863E+3   1.601227E+2   1.601227E+2   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   1.233973E-1   -1.400810E-1   1.675232E-4   3.125290E-7   -3.125290E-7   1.675232E-4   1.675235E-4   1.068901E-1   9.010689E+1   
2.509555E+3   1.600275E+2   1.600275E+2   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   1.244407E-1   -1.403482E-1   1.683423E-4   -2.845002E-7   2.845002E-7   1.683423E-4   1.683426E-4   -9.683033E-2   8.990317E+1   
2.531191E+3   1.601081E+2   1.601081E+2   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   1.255620E-1   -1.413697E-1   1.697009E-4   -4.460780E-7   4.460780E-7   1.697009E-4   1.697015E-4   -1.506081E-1   8.984939E+1   
2.552917E+3   1.600074E+2   1.600074E+2   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   1.257788E-1   -1.437177E-1   1.713641E-4   9.286752E-7   -9.286752E-7   1.713641E-4   1.713666E-4   3.105005E-1   9.031050E+1   
2.574570E+3   1.600363E+2   1.600363E+2   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   1.278306E-1   -1.455676E-1   1.738375E-4   6.205388E-7   -6.205388E-7   1.738375E-4   1.738386E-4   2.045249E-1   9.020452E+1   
2.596287E+3   1.600543E+2   1.600543E+2   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   1.283173E-1   -1.469226E-1   1.750209E-4   1.146363E-6   -1.146363E-6   1.750209E-4   1.750247E-4   3.752742E-1   9.037527E+1   
2.617997E+3   1.600001E+2   1.600001E+2   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   1.285089E-1   -1.478934E-1   1.757716E-4   1.639380E-6   -1.639380E-6   1.757716E-4   1.757793E-4   5.343685E-1   9.053437E+1   
2.640165E+3   1.599932E+2   1.599932E+2   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   1.299591E-1   -1.489835E-1   1.773782E-4   1.279388E-6   -1.279388E-6   1.773782E-4   1.773828E-4   4.132540E-1   9.041325E+1   
2.661906E+3   1.600167E+2   1.600167E+2   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.490000E+2   -6.490000E+2   1.302575E-1   -1.503888E-1   1.784779E-4   1.977436E-6   -1.977436E-6   1.784779E-4   1.784888E-4   6.347794E-1   9.063478E+1   
2.683594E+3   1.600299E+2   1.600299E+2   -7.000000E+2   -7.000000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   1.319528E-1   -1.519680E-1   1.805545E-4   1.755954E-6   -1.755954E-6   1.805545E-4   1.805631E-4   5.572034E-1   9.055720E+1   
2.705272E+3   1.599911E+2   1.599911E+2   -7.500000E+2   -7.500000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   1.338595E-1   -1.541288E-1   1.831407E-4   1.758414E-6   -1.758414E-6   1.831407E-4   1.831492E-4   5.501049E-1   9.055010E+1   
2.726990E+3   1.600380E+2   1.600380E+2   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   1.334691E-1   -1.555260E-1   1.838093E-4   2.960574E-6   -2.960574E-6   1.838093E-4   1.838331E-4   9.227702E-1   9.092277E+1   
2.748697E+3   1.600960E+2   1.600960E+2   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   1.348736E-1   -1.569219E-1   1.855867E-4   2.834379E-6   -2.834379E-6   1.855867E-4   1.856084E-4   8.749833E-1   9.087498E+1   
2.770349E+3   1.600107E+2   1.600107E+2   -9.000000E+2   -9.000000E+2   9.000000E+1   -9.000000E+2   -9.000000E+2   1.349945E-1   -1.583399E-1   1.865850E-4   3.672013E-6   -3.672013E-6   1.865850E-4   1.866211E-4   1.127442E+0   9.112744E+1   
2.792072E+3   1.599958E+2   1.599958E+2   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.490000E+2   -9.490000E+2   1.352632E-1   -1.600641E-1   1.878741E-4   4.600459E-6   -4.600459E-6   1.878741E-4   1.879304E-4   1.402717E+0   9.140272E+1   
2.813746E+3   1.600844E+2   1.600844E+2   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   1.360799E-1   -1.612027E-1   1.891206E-4   4.740832E-6   -4.740832E-6   1.891206E-4   1.891800E-4   1.435977E+0   9.143598E+1   
2.835619E+3   1.600497E+2   1.600497E+2   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   1.373441E-1   -1.624175E-1   1.906933E-4   4.600011E-6   -4.600011E-6   1.906933E-4   1.907488E-4   1.381853E+0   9.138185E+1   
2.857459E+3   1.600117E+2   1.600117E+2   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.100000E+3   -1.100000E+3   1.393388E-1   -1.650908E-1   1.936677E-4   4.872400E-6   -4.872400E-6   1.936677E-4   1.937290E-4   1.441175E+0   9.144118E+1   
2.879332E+3   1.600547E+2   1.600547E+2   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   1.385384E-1   -1.655877E-1   1.934965E-4   5.789248E-6   -5.789248E-6   1.934965E-4   1.935830E-4   1.713729E+0   9.171373E+1   
2.901713E+3   1.601065E+2   1.601065E+2   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   1.404074E-1   -1.672712E-1   1.957484E-4   5.507523E-6   -5.507523E-6   1.957484E-4   1.958259E-4   1.611633E+0   9.161163E+1   
2.923556E+3   1.600568E+2   1.600568E+2   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   1.418578E-1   -1.686938E-1   1.975716E-4   5.364847E-6   -5.364847E-6   1.975716E-4   1.976444E-4   1.555424E+0   9.155542E+1   
2.945350E+3   1.600573E+2   1.600573E+2   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   1.424672E-1   -1.713287E-1   1.996644E-4   6.636707E-6   -6.636707E-6   1.996644E-4   1.997747E-4   1.903771E+0   9.190377E+1   
2.967681E+3   1.600193E+2   1.600193E+2   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   1.444661E-1   -1.729678E-1   2.019678E-4   6.229808E-6   -6.229808E-6   2.019678E-4   2.020638E-4   1.766760E+0   9.176676E+1   
2.989747E+3   1.600769E+2   1.600769E+2   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   1.438982E-1   -1.732963E-1   2.018307E-4   6.864650E-6   -6.864650E-6   2.018307E-4   2.019474E-4   1.947989E+0   9.194799E+1   
3.011621E+3   1.599683E+2   1.599683E+2   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   1.454641E-1   -1.747085E-1   2.037185E-4   6.629710E-6   -6.629710E-6   2.037185E-4   2.038264E-4   1.863946E+0   9.186395E+1   
3.034464E+3   1.600422E+2   1.600422E+2   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   1.458317E-1   -1.768218E-1   2.053221E-4   7.739509E-6   -7.739509E-6   2.053221E-4   2.054680E-4   2.158712E+0   9.215871E+1   
3.056538E+3   1.600025E+2   1.600025E+2   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   1.470923E-1   -1.777536E-1   2.067083E-4   7.416261E-6   -7.416261E-6   2.067083E-4   2.068413E-4   2.054771E+0   9.205477E+1   
3.078660E+3   1.600220E+2   1.600220E+2   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   1.470823E-1   -1.793934E-1   2.077702E-4   8.495681E-6   -8.495681E-6   2.077702E-4   2.079438E-4   2.341509E+0   9.234151E+1   
3.101998E+3   1.600684E+2   1.600684E+2   -1.650000E+3   -1.650000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   1.486043E-1   -1.804909E-1   2.094259E-4   8.087535E-6   -8.087535E-6   2.094259E-4   2.095820E-4   2.211529E+0   9.221153E+1   
3.124148E+3   1.600741E+2   1.600741E+2   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   1.496462E-1   -1.839856E-1   2.123462E-4   9.601664E-6   -9.601664E-6   2.123462E-4   2.125631E-4   2.588982E+0   9.258898E+1   
3.146279E+3   1.600382E+2   1.600382E+2   -1.750000E+3   -1.750000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   1.502280E-1   -1.845882E-1   2.130983E-4   9.565256E-6   -9.565256E-6   2.130983E-4   2.133129E-4   2.570087E+0   9.257009E+1   
3.169402E+3   1.600573E+2   1.600573E+2   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.798000E+3   -1.798000E+3   1.511556E-1   -1.854713E-1   2.142470E-4   9.456575E-6   -9.456575E-6   2.142470E-4   2.144556E-4   2.527319E+0   9.252732E+1   
3.191978E+3   1.600372E+2   1.600372E+2   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.848000E+3   -1.848000E+3   1.532933E-1   -1.877258E-1   2.170369E-4   9.349346E-6   -9.349346E-6   2.170369E-4   2.172382E-4   2.466618E+0   9.246662E+1   
3.214503E+3   1.600424E+2   1.600424E+2   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   1.546657E-1   -1.892423E-1   2.188731E-4   9.325686E-6   -9.325686E-6   2.188731E-4   2.190717E-4   2.439768E+0   9.243977E+1   
3.237355E+3   1.600049E+2   1.600049E+2   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   1.545057E-1   -1.911186E-1   2.199962E-4   1.067068E-5   -1.067068E-5   2.199962E-4   2.202548E-4   2.776895E+0   9.277689E+1   
3.259727E+3   1.599661E+2   1.599661E+2   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   1.557228E-1   -1.908145E-1   2.205506E-4   9.571706E-6   -9.571706E-6   2.205506E-4   2.207582E-4   2.485028E+0   9.248503E+1   
3.296798E+3   1.599548E+2   1.599548E+2   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.633243E-1   -2.073779E-1   2.360378E-4   1.477803E-5   -1.477803E-5   2.360378E-4   2.364999E-4   3.582542E+0   9.358254E+1   
3.322936E+3   1.600673E+2   1.600673E+2   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.734088E-1   -2.235109E-1   2.527797E-4   1.786657E-5   -1.786657E-5   2.527797E-4   2.534103E-4   4.042967E+0   9.404297E+1   
3.348556E+3   1.600755E+2   1.600755E+2   -3.499000E+3   -3.499000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.788847E-1   -2.371219E-1   2.650299E-4   2.271489E-5   -2.271489E-5   2.650299E-4   2.660015E-4   4.898674E+0   9.489867E+1   
3.375193E+3   1.599786E+2   1.599786E+2   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   1.803082E-1   -2.423688E-1   2.693272E-4   2.509230E-5   -2.509230E-5   2.693272E-4   2.704935E-4   5.322689E+0   9.532269E+1   
3.401311E+3   1.600003E+2   1.600003E+2   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   1.703672E-1   -2.364066E-1   2.592981E-4   2.854704E-5   -2.854704E-5   2.592981E-4   2.608648E-4   6.282593E+0   9.628259E+1   
3.426037E+3   1.599808E+2   1.599808E+2   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   1.543907E-1   -2.204049E-1   2.389989E-4   2.990235E-5   -2.990235E-5   2.389989E-4   2.408623E-4   7.131504E+0   9.713150E+1   
3.451199E+3   1.600279E+2   1.600279E+2   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   1.381031E-1   -2.036546E-1   2.180199E-4   3.099831E-5   -3.099831E-5   2.180199E-4   2.202125E-4   8.092139E+0   9.809214E+1   
3.476907E+3   1.600760E+2   1.600760E+2   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   1.260348E-1   -1.923106E-1   2.031704E-4   3.250798E-5   -3.250798E-5   2.031704E-4   2.057547E-4   9.090472E+0   9.909047E+1   
3.501659E+3   1.600061E+2   1.600061E+2   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.214893E-1   -1.928852E-1   2.007345E-4   3.624559E-5   -3.624559E-5   2.007345E-4   2.039806E-4   1.023532E+1   1.002353E+2   
3.526400E+3   1.600464E+2   1.600464E+2   -7.001000E+3   -7.001000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.227389E-1   -1.975682E-1   2.045570E-4   3.838297E-5   -3.838297E-5   2.045570E-4   2.081269E-4   1.062738E+1   1.006274E+2   
3.551598E+3   1.600369E+2   1.600369E+2   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.301268E-1   -2.109130E-1   2.178159E-4   4.164317E-5   -4.164317E-5   2.178159E-4   2.217609E-4   1.082349E+1   1.008235E+2   
3.577257E+3   1.599985E+2   1.599985E+2   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.373159E-1   -2.240625E-1   2.308246E-4   4.492265E-5   -4.492265E-5   2.308246E-4   2.351553E-4   1.101313E+1   1.010131E+2   
3.602408E+3   1.600816E+2   1.600816E+2   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.455815E-1   -2.368309E-1   2.442507E-4   4.715677E-5   -4.715677E-5   2.442507E-4   2.487613E-4   1.092748E+1   1.009275E+2   
3.628120E+3   1.599997E+2   1.599997E+2   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.530307E-1   -2.528329E-1   2.592781E-4   5.210875E-5   -5.210875E-5   2.592781E-4   2.644626E-4   1.136371E+1   1.013637E+2   
3.653833E+3   1.599757E+2   1.599757E+2   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.642133E-1   -2.698716E-1   2.772888E-4   5.497716E-5   -5.497716E-5   2.772888E-4   2.826863E-4   1.121441E+1   1.012144E+2   
3.679074E+3   1.600114E+2   1.600114E+2   -1.000000E+4   -1.000000E+4   9.000000E+1   -9.999000E+3   -9.999000E+3   1.785012E-1   -2.909169E-1   2.998289E-4   5.816819E-5   -5.816819E-5   2.998289E-4   3.054192E-4   1.097926E+1   1.009793E+2   
3.715593E+3   1.600977E+2   1.600977E+2   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.660411E-1   -2.711550E-1   2.792548E-4   5.446432E-5   -5.446432E-5   2.792548E-4   2.845164E-4   1.103611E+1   1.010361E+2   
3.739806E+3   1.600473E+2   1.600473E+2   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.577062E-1   -2.532178E-1   2.624194E-4   4.890224E-5   -4.890224E-5   2.624194E-4   2.669370E-4   1.055607E+1   1.005561E+2   
3.764532E+3   1.600589E+2   1.600589E+2   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.463488E-1   -2.357534E-1   2.440234E-4   4.588484E-5   -4.588484E-5   2.440234E-4   2.482999E-4   1.064925E+1   1.006492E+2   
3.789187E+3   1.600177E+2   1.600177E+2   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.288269E-1   -2.134561E-1   2.186685E-4   4.426715E-5   -4.426715E-5   2.186685E-4   2.231042E-4   1.144427E+1   1.014443E+2   
3.813940E+3   1.600625E+2   1.600625E+2   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.200735E-1   -2.008717E-1   2.050607E-4   4.251417E-5   -4.251417E-5   2.050607E-4   2.094214E-4   1.171290E+1   1.017129E+2   
3.839143E+3   1.600683E+2   1.600683E+2   -7.000000E+3   -7.000000E+3   9.000000E+1   -6.999000E+3   -6.999000E+3   1.103160E-1   -1.824699E-1   1.870432E-4   3.770056E-5   -3.770056E-5   1.870432E-4   1.908048E-4   1.139589E+1   1.013959E+2   
3.863835E+3   1.600603E+2   1.600603E+2   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.022442E-1   -1.675478E-1   1.723343E-4   3.391500E-5   -3.391500E-5   1.723343E-4   1.756398E-4   1.113341E+1   1.011334E+2   
3.887964E+3   1.600341E+2   1.600341E+2   -5.999000E+3   -5.999000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   8.980323E-2   -1.484987E-1   1.522362E-4   3.066303E-5   -3.066303E-5   1.522362E-4   1.552936E-4   1.138800E+1   1.013880E+2   
3.912712E+3   1.600403E+2   1.600403E+2   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   7.843493E-2   -1.316942E-1   1.342632E-4   2.808503E-5   -2.808503E-5   1.342632E-4   1.371691E-4   1.181472E+1   1.018147E+2   
3.937355E+3   1.600163E+2   1.600163E+2   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   6.893203E-2   -1.161456E-1   1.182614E-4   2.494846E-5   -2.494846E-5   1.182614E-4   1.208643E-4   1.191246E+1   1.019125E+2   
3.962098E+3   1.600188E+2   1.600188E+2   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   5.923557E-2   -9.806845E-2   1.004931E-4   2.030192E-5   -2.030192E-5   1.004931E-4   1.025234E-4   1.142134E+1   1.014213E+2   
3.986800E+3   1.600048E+2   1.600048E+2   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.999000E+3   -3.999000E+3   4.540216E-2   -7.986765E-2   8.008669E-5   1.863436E-5   -1.863436E-5   8.008669E-5   8.222602E-5   1.309838E+1   1.030984E+2   
4.011562E+3   1.599609E+2   1.599609E+2   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   3.473953E-2   -6.344077E-2   6.279590E-5   1.578135E-5   -1.578135E-5   6.279590E-5   6.474856E-5   1.410696E+1   1.041070E+2   
4.035755E+3   1.600569E+2   1.600569E+2   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   2.431224E-2   -4.471248E-2   4.415173E-5   1.124967E-5   -1.124967E-5   4.415173E-5   4.556238E-5   1.429456E+1   1.042946E+2   
4.060450E+3   1.600183E+2   1.600183E+2   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.239848E-2   -2.841254E-2   2.617010E-5   9.405015E-6   -9.405015E-6   2.617010E-5   2.780878E-5   1.976743E+1   1.097674E+2   
4.085094E+3   1.600984E+2   1.600984E+2   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   4.192651E-3   -1.199412E-2   1.040374E-5   4.740404E-6   -4.740404E-6   1.040374E-5   1.143281E-5   2.449611E+1   1.144961E+2   
4.118794E+3   1.599929E+2   1.599929E+2   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   2.324581E-3   -9.508170E-3   7.629735E-6   4.496841E-6   -4.496841E-6   7.629735E-6   8.856322E-6   3.051440E+1   1.205144E+2   
4.140878E+3   1.600433E+2   1.600433E+2   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.899000E+3   -1.899000E+3   3.421062E-3   -8.631044E-3   7.736368E-6   3.112409E-6   -3.112409E-6   7.736368E-6   8.338973E-6   2.191536E+1   1.119154E+2   
4.162997E+3   1.599123E+2   1.599123E+2   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.849000E+3   -1.849000E+3   1.545323E-3   -5.445905E-3   4.502251E-6   2.417410E-6   -2.417410E-6   4.502251E-6   5.110199E-6   2.823284E+1   1.182328E+2   
4.184729E+3   1.600146E+2   1.600146E+2   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.798000E+3   -1.798000E+3   6.783220E-4   -3.999677E-3   3.024317E-6   2.113168E-6   -2.113168E-6   3.024317E-6   3.689441E-6   3.494298E+1   1.249430E+2   
4.206757E+3   1.599900E+2   1.599900E+2   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   -1.395903E-4   -2.100008E-3   1.281411E-6   1.476171E-6   -1.476171E-6   1.281411E-6   1.954763E-6   4.903992E+1   1.390399E+2   
4.228843E+3   1.600553E+2   1.600553E+2   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   -2.048465E-3   7.123767E-4   -1.730421E-6   1.049377E-6   -1.049377E-6   -1.730421E-6   2.023746E-6   1.487662E+2   2.387662E+2   
4.250724E+3   1.600301E+2   1.600301E+2   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   -2.705618E-3   8.670010E-4   -2.237408E-6   1.434339E-6   -1.434339E-6   -2.237408E-6   2.657691E-6   1.473372E+2   2.373372E+2   
4.272606E+3   1.600711E+2   1.600711E+2   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.599000E+3   -1.599000E+3   -4.057968E-3   1.356951E-3   -3.392593E-6   2.114263E-6   -2.114263E-6   -3.392593E-6   3.997474E-6   1.480689E+2   2.380689E+2   
4.294701E+3   1.600203E+2   1.600203E+2   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   -7.887987E-3   4.665422E-3   -7.915262E-6   2.784079E-6   -2.784079E-6   -7.915262E-6   8.390618E-6   1.606214E+2   2.506214E+2   
4.316573E+3   1.600307E+2   1.600307E+2   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   -5.123463E-3   7.104741E-3   -7.794807E-6   -8.554069E-7   8.554069E-7   -7.794807E-6   7.841603E-6   -1.737374E+2   -8.373739E+1   
4.338631E+3   1.600722E+2   1.600722E+2   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   -7.132352E-3   7.437919E-3   -9.253791E-6   4.126077E-7   -4.126077E-7   -9.253791E-6   9.262985E-6   1.774470E+2   2.674470E+2   
4.360666E+3   1.600719E+2   1.600719E+2   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   -8.040155E-3   9.759126E-3   -1.132682E-5   -4.334925E-7   4.334925E-7   -1.132682E-5   1.133511E-5   -1.778083E+2   -8.780828E+1   
4.382438E+3   1.599769E+2   1.599769E+2   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   -8.682584E-3   1.053470E-2   -1.222912E-5   -4.653805E-7   4.653805E-7   -1.222912E-5   1.223797E-5   -1.778207E+2   -8.782065E+1   
4.404561E+3   1.600191E+2   1.600191E+2   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   -9.354466E-3   1.331027E-2   -1.445221E-5   -1.783028E-6   1.783028E-6   -1.445221E-5   1.456178E-5   -1.729667E+2   -8.296673E+1   
4.426709E+3   1.600196E+2   1.600196E+2   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   -1.316884E-2   1.462887E-2   -1.766922E-5   1.761407E-7   -1.761407E-7   -1.766922E-5   1.767010E-5   1.794288E+2   2.694288E+2   
4.448791E+3   1.599944E+2   1.599944E+2   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   -1.159468E-2   1.548329E-2   -1.725248E-5   -1.546755E-6   1.546755E-6   -1.725248E-5   1.732167E-5   -1.748769E+2   -8.487690E+1   
4.470937E+3   1.599842E+2   1.599842E+2   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   -1.359590E-2   1.773976E-2   -1.995933E-5   -1.541803E-6   1.541803E-6   -1.995933E-5   2.001880E-5   -1.755828E+2   -8.558283E+1   
4.493000E+3   1.601142E+2   1.601142E+2   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.100000E+3   -1.100000E+3   -1.428527E-2   2.045304E-2   -2.215267E-5   -2.805793E-6   2.805793E-6   -2.215267E-5   2.232965E-5   -1.727815E+2   -8.278152E+1   
4.515032E+3   1.600233E+2   1.600233E+2   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.050000E+3   -1.050000E+3   -1.499610E-2   2.147283E-2   -2.325632E-5   -2.946748E-6   2.946748E-6   -2.325632E-5   2.344226E-5   -1.727787E+2   -8.277868E+1   
4.537097E+3   1.599811E+2   1.599811E+2   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   -1.543727E-2   2.308781E-2   -2.458089E-5   -3.676269E-6   3.676269E-6   -2.458089E-5   2.485428E-5   -1.714940E+2   -8.149400E+1   
4.559051E+3   1.600798E+2   1.600798E+2   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   -1.637575E-2   2.432941E-2   -2.596974E-5   -3.793864E-6   3.793864E-6   -2.596974E-5   2.624540E-5   -1.716886E+2   -8.168858E+1   
4.580748E+3   1.600363E+2   1.600363E+2   -9.000000E+2   -9.000000E+2   9.000000E+1   -8.990000E+2   -8.990000E+2   -1.744493E-2   2.544553E-2   -2.735768E-5   -3.732759E-6   3.732759E-6   -2.735768E-5   2.761116E-5   -1.722304E+2   -8.223038E+1   
4.602593E+3   1.599868E+2   1.599868E+2   -8.510000E+2   -8.510000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   -1.868744E-2   2.786738E-2   -2.970318E-5   -4.397095E-6   4.397095E-6   -2.970318E-5   3.002687E-5   -1.715794E+2   -8.157940E+1   
4.624222E+3   1.599597E+2   1.599597E+2   -8.000000E+2   -8.000000E+2   9.000000E+1   -8.000000E+2   -8.000000E+2   -1.889545E-2   2.948356E-2   -3.088438E-5   -5.299854E-6   5.299854E-6   -3.088438E-5   3.133581E-5   -1.702627E+2   -8.026271E+1   
4.645948E+3   1.600399E+2   1.600399E+2   -7.510000E+2   -7.510000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   -1.957346E-2   3.033430E-2   -3.185764E-5   -5.354571E-6   5.354571E-6   -3.185764E-5   3.230450E-5   -1.704590E+2   -8.045901E+1   
4.667821E+3   1.600488E+2   1.600488E+2   -7.010000E+2   -7.010000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   -2.134336E-2   3.145470E-2   -3.368158E-5   -4.777977E-6   4.777977E-6   -3.368158E-5   3.401878E-5   -1.719260E+2   -8.192605E+1   
4.689801E+3   1.600241E+2   1.600241E+2   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.500000E+2   -6.500000E+2   -2.334091E-2   3.307948E-2   -3.597476E-5   -4.362765E-6   4.362765E-6   -3.597476E-5   3.623834E-5   -1.730853E+2   -8.308534E+1   
4.711484E+3   1.600346E+2   1.600346E+2   -6.000000E+2   -6.000000E+2   9.000000E+1   -6.000000E+2   -6.000000E+2   -2.396831E-2   3.622594E-2   -3.841190E-5   -5.955788E-6   5.955788E-6   -3.841190E-5   3.887088E-5   -1.711864E+2   -8.118644E+1   
4.733115E+3   1.600266E+2   1.600266E+2   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   -2.438434E-2   3.631523E-2   -3.872726E-5   -5.706455E-6   5.706455E-6   -3.872726E-5   3.914542E-5   -1.716178E+2   -8.161779E+1   
4.754796E+3   1.600052E+2   1.600052E+2   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   -2.507646E-2   3.926257E-2   -4.107473E-5   -7.121433E-6   7.121433E-6   -4.107473E-5   4.168751E-5   -1.701640E+2   -8.016398E+1   
4.776437E+3   1.600720E+2   1.600720E+2   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   -2.733110E-2   4.035199E-2   -4.317818E-5   -6.166061E-6   6.166061E-6   -4.317818E-5   4.361623E-5   -1.718728E+2   -8.187283E+1   
4.798121E+3   1.599846E+2   1.599846E+2   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   -2.739459E-2   4.131442E-2   -4.384426E-5   -6.748310E-6   6.748310E-6   -4.384426E-5   4.436056E-5   -1.712500E+2   -8.124996E+1   
4.819796E+3   1.600177E+2   1.600177E+2   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   -2.756732E-2   4.338068E-2   -4.529679E-5   -7.971417E-6   7.971417E-6   -4.529679E-5   4.599285E-5   -1.700192E+2   -8.001917E+1   
4.841495E+3   1.600174E+2   1.600174E+2   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   -2.881044E-2   4.450384E-2   -4.679684E-5   -7.786256E-6   7.786256E-6   -4.679684E-5   4.744018E-5   -1.705534E+2   -8.055343E+1   
4.863222E+3   1.600949E+2   1.600949E+2   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   -3.062422E-2   4.583902E-2   -4.878779E-5   -7.317634E-6   7.317634E-6   -4.878779E-5   4.933352E-5   -1.714698E+2   -8.146985E+1   
4.884950E+3   1.600073E+2   1.600073E+2   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   -3.135253E-2   4.705149E-2   -5.002774E-5   -7.571631E-6   7.571631E-6   -5.002774E-5   5.059747E-5   -1.713937E+2   -8.139368E+1   
4.906579E+3   1.600669E+2   1.600669E+2   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   -3.306078E-2   4.870395E-2   -5.216009E-5   -7.388493E-6   7.388493E-6   -5.216009E-5   5.268078E-5   -1.719377E+2   -8.193767E+1   
4.928264E+3   1.600023E+2   1.600023E+2   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   -3.309972E-2   4.999986E-2   -5.302817E-5   -8.206916E-6   8.206916E-6   -5.302817E-5   5.365948E-5   -1.712024E+2   -8.120240E+1   
4.949862E+3   1.600040E+2   1.600040E+2   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   -3.395905E-2   5.165438E-2   -5.463702E-5   -8.653010E-6   8.653010E-6   -5.463702E-5   5.531798E-5   -1.710007E+2   -8.100066E+1   
4.982899E+3   1.600123E+2   1.600123E+2   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.600000E+1   -4.600000E+1   -3.458490E-2   5.188051E-2   -5.517123E-5   -8.337949E-6   8.337949E-6   -5.517123E-5   5.579772E-5   -1.714060E+2   -8.140600E+1   
5.005190E+3   1.601056E+2   1.601056E+2   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   -3.359490E-2   5.309787E-2   -5.535202E-5   -9.866053E-6   9.866053E-6   -5.535202E-5   5.622441E-5   -1.698936E+2   -7.989362E+1   
5.027495E+3   1.599808E+2   1.599808E+2   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   -3.428702E-2   5.367925E-2   -5.615856E-5   -9.734232E-6   9.734232E-6   -5.615856E-5   5.699596E-5   -1.701664E+2   -8.016636E+1   
5.049761E+3   1.601280E+2   1.601280E+2   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   -3.365533E-2   5.294478E-2   -5.528967E-5   -9.721276E-6   9.721276E-6   -5.528967E-5   5.613778E-5   -1.700279E+2   -8.002793E+1   
5.071921E+3   1.599817E+2   1.599817E+2   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   -3.310617E-2   5.290091E-2   -5.492158E-5   -1.009877E-5   1.009877E-5   -5.492158E-5   5.584233E-5   -1.695811E+2   -7.958105E+1   
5.094198E+3   1.600404E+2   1.600404E+2   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   -3.363508E-2   5.265119E-2   -5.508594E-5   -9.544315E-6   9.544315E-6   -5.508594E-5   5.590666E-5   -1.701704E+2   -8.017039E+1   
5.116449E+3   1.600233E+2   1.600233E+2   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   -3.342369E-2   5.192131E-2   -5.447989E-5   -9.223487E-6   9.223487E-6   -5.447989E-5   5.525514E-5   -1.703909E+2   -8.039090E+1   
5.138735E+3   1.600899E+2   1.600899E+2   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   -3.338043E-2   5.402099E-2   -5.582064E-5   -1.062819E-5   1.062819E-5   -5.582064E-5   5.682343E-5   -1.692200E+2   -7.921997E+1   
5.161030E+3   1.600505E+2   1.600505E+2   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   -3.372005E-2   5.301073E-2   -5.537264E-5   -9.716526E-6   9.716526E-6   -5.537264E-5   5.621868E-5   -1.700473E+2   -8.004734E+1   
5.183216E+3   1.599594E+2   1.599594E+2   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   -3.450698E-2   5.291838E-2   -5.579901E-5   -9.074112E-6   9.074112E-6   -5.579901E-5   5.653202E-5   -1.707633E+2   -8.076334E+1   
5.205472E+3   1.599954E+2   1.599954E+2   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   -3.412319E-2   5.279995E-2   -5.548460E-5   -9.280550E-6   9.280550E-6   -5.548460E-5   5.625539E-5   -1.705044E+2   -8.050441E+1   
5.227788E+3   1.599997E+2   1.599997E+2   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   -3.473983E-2   5.299693E-2   -5.599412E-5   -8.953242E-6   8.953242E-6   -5.599412E-5   5.670540E-5   -1.709155E+2   -8.091553E+1   
5.250031E+3   1.600473E+2   1.600473E+2   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   -3.339886E-2   5.324053E-2   -5.532373E-5   -1.010432E-5   1.010432E-5   -5.532373E-5   5.623889E-5   -1.696496E+2   -7.964958E+1   
5.272269E+3   1.600203E+2   1.600203E+2   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   -3.488249E-2   5.347338E-2   -5.639263E-5   -9.159214E-6   9.159214E-6   -5.639263E-5   5.713160E-5   -1.707747E+2   -8.077466E+1   
5.294451E+3   1.599823E+2   1.599823E+2   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   -3.360532E-2   5.274904E-2   -5.513127E-5   -9.630292E-6   9.630292E-6   -5.513127E-5   5.596606E-5   -1.700916E+2   -8.009158E+1   
5.316700E+3   1.599619E+2   1.599619E+2   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   -3.449288E-2   5.304754E-2   -5.587441E-5   -9.168982E-6   9.168982E-6   -5.587441E-5   5.662173E-5   -1.706808E+2   -8.068083E+1   
5.338873E+3   1.599554E+2   1.599554E+2   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   -3.465147E-2   5.475516E-2   -5.708461E-5   -1.016808E-5   1.016808E-5   -5.708461E-5   5.798312E-5   -1.699002E+2   -7.990024E+1   
5.361114E+3   1.600285E+2   1.600285E+2   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   -3.415815E-2   5.355683E-2   -5.599916E-5   -9.749518E-6   9.749518E-6   -5.599916E-5   5.684153E-5   -1.701237E+2   -8.012373E+1   
5.383385E+3   1.599499E+2   1.599499E+2   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   -3.430696E-2   5.445480E-2   -5.667600E-5   -1.022652E-5   1.022652E-5   -5.667600E-5   5.759124E-5   -1.697717E+2   -7.977171E+1   
5.405530E+3   1.600579E+2   1.600579E+2   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   -3.521721E-2   5.509416E-2   -5.765517E-5   -9.971269E-6   9.971269E-6   -5.765517E-5   5.851106E-5   -1.701879E+2   -8.018795E+1   
5.427657E+3   1.600243E+2   1.600243E+2   -7.000000E+0   -7.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   -3.402194E-2   5.456402E-2   -5.657093E-5   -1.050873E-5   1.050873E-5   -5.657093E-5   5.753871E-5   -1.694766E+2   -7.947657E+1   
5.448733E+3   1.600057E+2   1.600057E+2   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   -3.338136E-2   5.358998E-2   -5.554050E-5   -1.034572E-5   1.034572E-5   -5.554050E-5   5.649585E-5   -1.694482E+2   -7.944825E+1   
5.470804E+3   1.599802E+2   1.599802E+2   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   -3.480089E-2   5.422871E-2   -5.683412E-5   -9.713375E-6   9.713375E-6   -5.683412E-5   5.765819E-5   -1.703014E+2   -8.030143E+1   
5.492848E+3   1.600678E+2   1.600678E+2   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   -3.564120E-2   5.373048E-2   -5.702915E-5   -8.766131E-6   8.766131E-6   -5.702915E-5   5.769896E-5   -1.712613E+2   -8.126128E+1   
5.514898E+3   1.599389E+2   1.599389E+2   0.000000E+0   0.000000E+0   9.000000E+1   0.000000E+0   0.000000E+0   -3.539209E-2   5.350805E-2   -5.673027E-5   -8.804965E-6   8.804965E-6   -5.673027E-5   5.740950E-5   -1.711777E+2   -8.117766E+1   
5.536970E+3   1.600813E+2   1.600813E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   -3.504295E-2   5.470883E-2   -5.729647E-5   -9.848230E-6   9.848230E-6   -5.729647E-5   5.813668E-5   -1.702472E+2   -8.024719E+1   
5.558455E+3   1.600129E+2   1.600129E+2   3.000000E+0   3.000000E+0   9.000000E+1   3.000000E+0   3.000000E+0   -3.479905E-2   5.450636E-2   -5.701382E-5   -9.896255E-6   9.896255E-6   -5.701382E-5   5.786632E-5   -1.701529E+2   -8.015291E+1   
5.580186E+3   1.600324E+2   1.600324E+2   5.000000E+0   5.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   -3.445728E-2   5.392436E-2   -5.642347E-5   -9.768546E-6   9.768546E-6   -5.642347E-5   5.726283E-5   -1.701778E+2   -8.017779E+1   
5.601918E+3   1.600472E+2   1.600472E+2   7.000000E+0   7.000000E+0   9.000000E+1   8.000000E+0   8.000000E+0   -3.468431E-2   5.445973E-2   -5.691251E-5   -9.950635E-6   9.950635E-6   -5.691251E-5   5.777585E-5   -1.700826E+2   -8.008260E+1   
5.623703E+3   1.600407E+2   1.600407E+2   9.000000E+0   9.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   -3.483771E-2   5.417747E-2   -5.682352E-5   -9.652647E-6   9.652647E-6   -5.682352E-5   5.763754E-5   -1.703592E+2   -8.035916E+1   
5.645741E+3   1.600490E+2   1.600490E+2   1.100000E+1   1.100000E+1   9.000000E+1   1.100000E+1   1.100000E+1   -3.534667E-2   5.436338E-2   -5.725926E-5   -9.397744E-6   9.397744E-6   -5.725926E-5   5.802534E-5   -1.706794E+2   -8.067936E+1   
5.667777E+3   1.600365E+2   1.600365E+2   1.300000E+1   1.300000E+1   9.000000E+1   1.300000E+1   1.300000E+1   -3.484599E-2   5.440388E-2   -5.697609E-5   -9.794545E-6   9.794545E-6   -5.697609E-5   5.781184E-5   -1.702458E+2   -8.024584E+1   
5.689756E+3   1.600676E+2   1.600676E+2   1.500000E+1   1.500000E+1   9.000000E+1   1.500000E+1   1.500000E+1   -3.570256E-2   5.395228E-2   -5.721154E-5   -8.865752E-6   8.865752E-6   -5.721154E-5   5.789440E-5   -1.711913E+2   -8.119126E+1   
5.711778E+3   1.600772E+2   1.600772E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   -3.595044E-2   5.508466E-2   -5.810229E-5   -9.422734E-6   9.422734E-6   -5.810229E-5   5.886140E-5   -1.707883E+2   -8.078826E+1   
5.733613E+3   1.600590E+2   1.600590E+2   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   -3.450484E-2   5.604122E-2   -5.783156E-5   -1.111732E-5   1.111732E-5   -5.783156E-5   5.889044E-5   -1.691184E+2   -7.911843E+1   
5.755447E+3   1.600222E+2   1.600222E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   -3.647906E-2   5.487541E-2   -5.829283E-5   -8.894951E-6   8.894951E-6   -5.829283E-5   5.896757E-5   -1.713241E+2   -8.132411E+1   
5.777362E+3   1.600040E+2   1.600040E+2   2.300000E+1   2.300000E+1   9.000000E+1   2.300000E+1   2.300000E+1   -3.535526E-2   5.472601E-2   -5.750075E-5   -9.628469E-6   9.628469E-6   -5.750075E-5   5.830132E-5   -1.704940E+2   -8.049404E+1   
5.799395E+3   1.600252E+2   1.600252E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   -3.507455E-2   5.548473E-2   -5.782134E-5   -1.033212E-5   1.033212E-5   -5.782134E-5   5.873721E-5   -1.698687E+2   -7.986872E+1   
5.821331E+3   1.599767E+2   1.599767E+2   2.600000E+1   2.600000E+1   9.000000E+1   2.800000E+1   2.800000E+1   -3.606304E-2   5.468276E-2   -5.791016E-5   -9.076697E-6   9.076697E-6   -5.791016E-5   5.861717E-5   -1.710921E+2   -8.109207E+1   
5.843260E+3   1.600180E+2   1.600180E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   -3.564151E-2   5.658304E-2   -5.888718E-5   -1.063083E-5   1.063083E-5   -5.888718E-5   5.983907E-5   -1.697667E+2   -7.976669E+1   
5.865201E+3   1.600012E+2   1.600012E+2   3.000000E+1   3.000000E+1   9.000000E+1   3.100000E+1   3.100000E+1   -3.485981E-2   5.478951E-2   -5.723579E-5   -1.003644E-5   1.003644E-5   -5.723579E-5   5.810909E-5   -1.700542E+2   -8.005416E+1   
5.887143E+3   1.600167E+2   1.600167E+2   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   -3.634834E-2   5.582617E-2   -5.883124E-5   -9.613210E-6   9.613210E-6   -5.883124E-5   5.961148E-5   -1.707197E+2   -8.071970E+1   
5.909025E+3   1.600040E+2   1.600040E+2   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   -3.698954E-2   5.576265E-2   -5.918629E-5   -9.097434E-6   9.097434E-6   -5.918629E-5   5.988138E-5   -1.712615E+2   -8.126154E+1   
5.930900E+3   1.600116E+2   1.600116E+2   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   -3.503620E-2   5.557706E-2   -5.785777E-5   -1.042085E-5   1.042085E-5   -5.785777E-5   5.878874E-5   -1.697898E+2   -7.978984E+1   
5.952778E+3   1.600028E+2   1.600028E+2   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   -3.636523E-2   5.552612E-2   -5.864626E-5   -9.404558E-6   9.404558E-6   -5.864626E-5   5.939554E-5   -1.708896E+2   -8.088957E+1   
5.974623E+3   1.600181E+2   1.600181E+2   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   -3.787956E-2   5.460852E-2   -5.898486E-5   -7.684604E-6   7.684604E-6   -5.898486E-5   5.948334E-5   -1.725773E+2   -8.257726E+1   
5.996510E+3   1.600203E+2   1.600203E+2   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   -3.570655E-2   5.576235E-2   -5.839289E-5   -1.004618E-5   1.004618E-5   -5.839289E-5   5.925078E-5   -1.702381E+2   -8.023814E+1   
6.018326E+3   1.599749E+2   1.599749E+2   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   -3.635202E-2   5.648915E-2   -5.926531E-5   -1.004393E-5   1.004393E-5   -5.926531E-5   6.011038E-5   -1.703812E+2   -8.038125E+1   
6.040205E+3   1.599752E+2   1.599752E+2   4.600000E+1   4.600000E+1   9.000000E+1   4.700000E+1   4.700000E+1   -3.604464E-2   5.531687E-2   -5.831177E-5   -9.504874E-6   9.504874E-6   -5.831177E-5   5.908135E-5   -1.707422E+2   -8.074215E+1   
6.062129E+3   1.601019E+2   1.601019E+2   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   -3.623545E-2   5.664163E-2   -5.929254E-5   -1.022983E-5   1.022983E-5   -5.929254E-5   6.016856E-5   -1.702110E+2   -8.021104E+1   
6.096114E+3   1.600563E+2   1.600563E+2   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   -3.756632E-2   5.851458E-2   -6.133519E-5   -1.046996E-5   1.046996E-5   -6.133519E-5   6.222238E-5   -1.703129E+2   -8.031294E+1   
6.118752E+3   1.600586E+2   1.600586E+2   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   -3.692511E-2   5.789087E-2   -6.053254E-5   -1.053646E-5   1.053646E-5   -6.053254E-5   6.144270E-5   -1.701259E+2   -8.012587E+1   
6.140941E+3   1.600310E+2   1.600310E+2   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   -3.852107E-2   6.075848E-2   -6.338688E-5   -1.123080E-5   1.123080E-5   -6.338688E-5   6.437412E-5   -1.699527E+2   -7.995269E+1   
6.163270E+3   1.600423E+2   1.600423E+2   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   -3.864069E-2   6.303180E-2   -6.494143E-5   -1.262855E-5   1.262855E-5   -6.494143E-5   6.615791E-5   -1.689956E+2   -7.899556E+1   
6.186163E+3   1.600299E+2   1.600299E+2   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   -4.175650E-2   6.349783E-2   -6.717128E-5   -1.062868E-5   1.062868E-5   -6.717128E-5   6.800699E-5   -1.710085E+2   -8.100849E+1   
6.208478E+3   1.600016E+2   1.600016E+2   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   -4.228020E-2   6.512414E-2   -6.855426E-5   -1.130458E-5   1.130458E-5   -6.855426E-5   6.948007E-5   -1.706362E+2   -8.063621E+1   
6.230675E+3   1.600363E+2   1.600363E+2   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   -4.338773E-2   6.587547E-2   -6.972832E-5   -1.097661E-5   1.097661E-5   -6.972832E-5   7.058700E-5   -1.710539E+2   -8.105393E+1   
6.253287E+3   1.599468E+2   1.599468E+2   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   -4.282875E-2   6.804172E-2   -7.079359E-5   -1.280628E-5   1.280628E-5   -7.079359E-5   7.194257E-5   -1.697463E+2   -7.974630E+1   
6.275466E+3   1.599995E+2   1.599995E+2   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   -4.610319E-2   7.061266E-2   -7.449243E-5   -1.206521E-5   1.206521E-5   -7.449243E-5   7.546318E-5   -1.707999E+2   -8.079995E+1   
6.298076E+3   1.600072E+2   1.600072E+2   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   -4.551998E-2   7.044175E-2   -7.402055E-5   -1.238484E-5   1.238484E-5   -7.402055E-5   7.504949E-5   -1.705015E+2   -8.050147E+1   
6.321464E+3   1.600225E+2   1.600225E+2   5.980000E+2   5.980000E+2   9.000000E+1   5.990000E+2   5.990000E+2   -4.604335E-2   7.217392E-2   -7.547226E-5   -1.313017E-5   1.313017E-5   -7.547226E-5   7.660590E-5   -1.701308E+2   -8.013083E+1   
6.344091E+3   1.601399E+2   1.601399E+2   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   -4.674595E-2   7.255435E-2   -7.615441E-5   -1.285923E-5   1.285923E-5   -7.615441E-5   7.723246E-5   -1.704156E+2   -8.041560E+1   
6.366721E+3   1.600072E+2   1.600072E+2   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   -4.938717E-2   7.550906E-2   -7.971171E-5   -1.283741E-5   1.283741E-5   -7.971171E-5   8.073881E-5   -1.708512E+2   -8.085119E+1   
6.390095E+3   1.600066E+2   1.600066E+2   7.480000E+2   7.480000E+2   9.000000E+1   7.480000E+2   7.480000E+2   -4.901289E-2   7.716912E-2   -8.056149E-5   -1.419954E-5   1.419954E-5   -8.056149E-5   8.180331E-5   -1.700039E+2   -8.000388E+1   
6.412658E+3   1.600807E+2   1.600807E+2   7.970000E+2   7.970000E+2   9.000000E+1   7.980000E+2   7.980000E+2   -5.004710E-2   7.877364E-2   -8.224589E-5   -1.448359E-5   1.448359E-5   -8.224589E-5   8.351144E-5   -1.700126E+2   -8.001256E+1   
6.435291E+3   1.599839E+2   1.599839E+2   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   -5.159058E-2   8.066346E-2   -8.443097E-5   -1.457750E-5   1.457750E-5   -8.443097E-5   8.568017E-5   -1.702041E+2   -8.020413E+1   
6.458640E+3   1.600915E+2   1.600915E+2   8.970000E+2   8.970000E+2   9.000000E+1   8.980000E+2   8.980000E+2   -5.152371E-2   8.221093E-2   -8.539747E-5   -1.563865E-5   1.563865E-5   -8.539747E-5   8.681760E-5   -1.696225E+2   -7.962254E+1   
6.481322E+3   1.599574E+2   1.599574E+2   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   -5.279751E-2   8.261253E-2   -8.644656E-5   -1.495906E-5   1.495906E-5   -8.644656E-5   8.773130E-5   -1.701825E+2   -8.018253E+1   
6.503913E+3   1.600425E+2   1.600425E+2   9.980000E+2   9.980000E+2   9.000000E+1   9.980000E+2   9.980000E+2   -5.460760E-2   8.399678E-2   -8.846719E-5   -1.452525E-5   1.452525E-5   -8.846719E-5   8.965169E-5   -1.706759E+2   -8.067591E+1   
6.527365E+3   1.600565E+2   1.600565E+2   1.048000E+3   1.048000E+3   9.000000E+1   1.048000E+3   1.048000E+3   -5.606456E-2   8.651187E-2   -9.100600E-5   -1.509193E-5   1.509193E-5   -9.100600E-5   9.224889E-5   -1.705841E+2   -8.058408E+1   
6.550375E+3   1.599836E+2   1.599836E+2   1.097000E+3   1.097000E+3   9.000000E+1   1.098000E+3   1.098000E+3   -5.546662E-2   8.800318E-2   -9.160760E-5   -1.650916E-5   1.650916E-5   -9.160760E-5   9.308332E-5   -1.697840E+2   -7.978403E+1   
6.573439E+3   1.599430E+2   1.599430E+2   1.148000E+3   1.148000E+3   9.000000E+1   1.148000E+3   1.148000E+3   -5.696960E-2   8.852381E-2   -9.287589E-5   -1.573788E-5   1.573788E-5   -9.287589E-5   9.419985E-5   -1.703825E+2   -8.038255E+1   
6.597004E+3   1.600149E+2   1.600149E+2   1.198000E+3   1.198000E+3   9.000000E+1   1.198000E+3   1.198000E+3   -5.782124E-2   9.117699E-2   -9.513040E-5   -1.684256E-5   1.684256E-5   -9.513040E-5   9.660986E-5   -1.699600E+2   -7.995999E+1   
6.619839E+3   1.600393E+2   1.600393E+2   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   -5.770621E-2   9.330991E-2   -9.644844E-5   -1.832208E-5   1.832208E-5   -9.644844E-5   9.817331E-5   -1.692438E+2   -7.924382E+1   
6.642830E+3   1.600345E+2   1.600345E+2   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   -5.941688E-2   9.403734E-2   -9.797982E-5   -1.753239E-5   1.753239E-5   -9.797982E-5   9.953607E-5   -1.698549E+2   -7.985493E+1   
6.666377E+3   1.599596E+2   1.599596E+2   1.348000E+3   1.348000E+3   9.000000E+1   1.348000E+3   1.348000E+3   -6.052624E-2   9.639052E-2   -1.001983E-4   -1.825032E-5   1.825032E-5   -1.001983E-4   1.018468E-4   -1.696772E+2   -7.967719E+1   
6.688916E+3   1.600798E+2   1.600798E+2   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   -6.188810E-2   9.788224E-2   -1.020118E-4   -1.821828E-5   1.821828E-5   -1.020118E-4   1.036258E-4   -1.698743E+2   -7.987430E+1   
6.711432E+3   1.600024E+2   1.600024E+2   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   -6.321283E-2   9.962269E-2   -1.039643E-4   -1.837633E-5   1.837633E-5   -1.039643E-4   1.055759E-4   -1.699762E+2   -7.997615E+1   
6.734522E+3   1.600090E+2   1.600090E+2   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   -6.323307E-2   1.003424E-1   -1.044456E-4   -1.883190E-5   1.883190E-5   -1.044456E-4   1.061297E-4   -1.697792E+2   -7.977919E+1   
6.757075E+3   1.600703E+2   1.600703E+2   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   -6.584143E-2   1.025204E-1   -1.074767E-4   -1.832655E-5   1.832655E-5   -1.074767E-4   1.090280E-4   -1.703232E+2   -8.032319E+1   
6.779661E+3   1.600697E+2   1.600697E+2   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   -6.470997E-2   1.046786E-1   -1.081828E-4   -2.057444E-5   2.057444E-5   -1.081828E-4   1.101219E-4   -1.692320E+2   -7.923196E+1   
6.802723E+3   1.600145E+2   1.600145E+2   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   -6.648384E-2   1.056637E-1   -1.099211E-4   -1.990646E-5   1.990646E-5   -1.099211E-4   1.117091E-4   -1.697351E+2   -7.973512E+1   
6.825250E+3   1.600301E+2   1.600301E+2   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   -6.698698E-2   1.056874E-1   -1.102475E-4   -1.954977E-5   1.954977E-5   -1.102475E-4   1.119675E-4   -1.699445E+2   -7.994449E+1   
6.847791E+3   1.598789E+2   1.598789E+2   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   -6.767665E-2   1.087749E-1   -1.126848E-4   -2.105823E-5   2.105823E-5   -1.126848E-4   1.146356E-4   -1.694148E+2   -7.941482E+1   
6.870531E+3   1.599489E+2   1.599489E+2   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   -6.997239E-2   1.094039E-1   -1.145138E-4   -1.977141E-5   1.977141E-5   -1.145138E-4   1.162081E-4   -1.702042E+2   -8.020416E+1   
6.893117E+3   1.600442E+2   1.600442E+2   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   -7.049241E-2   1.121441E-1   -1.166200E-4   -2.117829E-5   2.117829E-5   -1.166200E-4   1.185274E-4   -1.697072E+2   -7.970721E+1   
6.915648E+3   1.600355E+2   1.600355E+2   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   -7.062707E-2   1.131090E-1   -1.173317E-4   -2.170950E-5   2.170950E-5   -1.173317E-4   1.193232E-4   -1.695173E+2   -7.951730E+1   
6.938524E+3   1.600603E+2   1.600603E+2   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   -7.224542E-2   1.142490E-1   -1.190747E-4   -2.125785E-5   2.125785E-5   -1.190747E-4   1.209573E-4   -1.698779E+2   -7.987789E+1   
6.961013E+3   1.599949E+2   1.599949E+2   1.999000E+3   1.999000E+3   9.000000E+1   2.000000E+3   2.000000E+3   -7.326335E-2   1.170592E-1   -1.215343E-4   -2.234218E-5   2.234218E-5   -1.215343E-4   1.235708E-4   -1.695834E+2   -7.958337E+1   
6.998974E+3   1.599751E+2   1.599751E+2   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   -8.210050E-2   1.303455E-1   -1.356510E-4   -2.449214E-5   2.449214E-5   -1.356510E-4   1.378444E-4   -1.697654E+2   -7.976536E+1   
7.025616E+3   1.599672E+2   1.599672E+2   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   -9.158044E-2   1.454756E-1   -1.513660E-4   -2.737211E-5   2.737211E-5   -1.513660E-4   1.538210E-4   -1.697498E+2   -7.974975E+1   
7.051516E+3   1.600703E+2   1.600703E+2   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -9.673389E-2   1.574141E-1   -1.623276E-4   -3.136553E-5   3.136553E-5   -1.623276E-4   1.653301E-4   -1.690639E+2   -7.906387E+1   
7.077358E+3   1.600229E+2   1.600229E+2   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -9.833077E-2   1.626677E-1   -1.667364E-4   -3.361902E-5   3.361902E-5   -1.667364E-4   1.700919E-4   -1.686003E+2   -7.860031E+1   
7.103883E+3   1.599731E+2   1.599731E+2   4.497000E+3   4.497000E+3   9.000000E+1   4.499000E+3   4.499000E+3   -8.727121E-2   1.544103E-1   -1.545210E-4   -3.640062E-5   3.640062E-5   -1.545210E-4   1.587505E-4   -1.667445E+2   -7.674446E+1   
7.129990E+3   1.599868E+2   1.599868E+2   4.997000E+3   4.997000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -7.066760E-2   1.379914E-1   -1.335624E-4   -3.794695E-5   3.794695E-5   -1.335624E-4   1.388484E-4   -1.641394E+2   -7.413940E+1   
7.155665E+3   1.600550E+2   1.600550E+2   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -5.683001E-2   1.252663E-1   -1.167196E-4   -3.986230E-5   3.986230E-5   -1.167196E-4   1.233388E-4   -1.611438E+2   -7.114383E+1   
7.182108E+3   1.600695E+2   1.600695E+2   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -4.630322E-2   1.162779E-1   -1.043574E-4   -4.177188E-5   4.177188E-5   -1.043574E-4   1.124071E-4   -1.581849E+2   -6.818490E+1   
7.208108E+3   1.600758E+2   1.600758E+2   6.497000E+3   6.497000E+3   9.000000E+1   6.499000E+3   6.499000E+3   -4.421607E-2   1.161226E-1   -1.029659E-4   -4.321411E-5   4.321411E-5   -1.029659E-4   1.116666E-4   -1.572325E+2   -6.723252E+1   
7.234265E+3   1.599941E+2   1.599941E+2   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -4.628972E-2   1.237084E-1   -1.091884E-4   -4.663973E-5   4.663973E-5   -1.091884E-4   1.187324E-4   -1.568703E+2   -6.687030E+1   
7.260198E+3   1.600181E+2   1.600181E+2   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -5.181392E-2   1.335926E-1   -1.190413E-4   -4.901591E-5   4.901591E-5   -1.190413E-4   1.287376E-4   -1.576203E+2   -6.762031E+1   
7.285591E+3   1.600584E+2   1.600584E+2   7.999000E+3   7.999000E+3   9.000000E+1   8.000000E+3   8.000000E+3   -5.984456E-2   1.458490E-1   -1.319886E-4   -5.108906E-5   5.108906E-5   -1.319886E-4   1.415312E-4   -1.588400E+2   -6.883999E+1   
7.312040E+3   1.600078E+2   1.600078E+2   8.497000E+3   8.497000E+3   9.000000E+1   8.499000E+3   8.499000E+3   -7.007210E-2   1.637948E-1   -1.499997E-4   -5.525692E-5   5.525692E-5   -1.499997E-4   1.598538E-4   -1.597772E+2   -6.977720E+1   
7.338436E+3   1.599510E+2   1.599510E+2   8.998000E+3   8.998000E+3   9.000000E+1   8.999000E+3   8.999000E+3   -7.654909E-2   1.782067E-1   -1.633904E-4   -5.988841E-5   5.988841E-5   -1.633904E-4   1.740202E-4   -1.598703E+2   -6.987031E+1   
7.364846E+3   1.600369E+2   1.600369E+2   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -8.968785E-2   1.985377E-1   -1.847547E-4   -6.346240E-5   6.346240E-5   -1.847547E-4   1.953504E-4   -1.610426E+2   -7.104264E+1   
7.390048E+3   1.600818E+2   1.600818E+2   9.999000E+3   9.999000E+3   9.000000E+1   1.000000E+4   1.000000E+4   -1.022298E-1   2.160577E-1   -2.039193E-4   -6.564003E-5   6.564003E-5   -2.039193E-4   2.142235E-4   -1.621570E+2   -7.215704E+1   
@@END Data.
@Time at end of measurement: 17:14:43
@Instrument  Changes:
@Emu Range: 20 uV
@END Instrument  Changes:
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -9499.000      -9999.000      250.000        Coercive Field: Field at which M//H changes sign
Ms  emu                                 2.998E-4       -2.039E-4      2.519E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -5.673E-5      1.596E-4       1.082E-4       Remanent Magnetization: M at H=0        
S                                       0.189          0.783          0.486          Squareness: Mr/Ms                       
S*                                      1.499          1.126          1.312          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
