@Filename: c:\vsm-lv\Will\data\AJA335e-FePtFeRh_1030nm_Tann_6\AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_130deg.VHD
@Measurement Controlfilename: C:\vsm-lv\Will\Recipes\10kOe OoP loop 130deg.VHC
@Signal Manipulation filename: c:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA335e-FePtFeRh_1030nm_Tann_6
@Date: 08 November 2019    (2019-08-11)
@Time: 15:32:54
@Test ID: AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_130deg
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 90.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Sample Temperature to 130.0530 [degC] and wait 60.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Applied Field to 9999.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 3:      Set Auto Range Signal to 12.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 5
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 5.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 10000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To: 50.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: 50.0000 [Oe] To: -50.0000 [Oe] Min Stepsize/Sweeprate =  2.0000 [Oe] Max Stepsize/Sweeprate =  2.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -50.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -10000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 4 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 20 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.706
@Y Coils Correction Factor: 0.964
@Sample Shape Correction Factor: 0.919
@Coil Angle Alpha: 42.300
@Coil Angle Beta: -47.320
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
15000.000000   1.000000
15249.000000   1.000524
15499.000000   1.000702
15750.000000   1.001233
16000.000000   1.001406
16250.000000   1.001585
16499.000000   1.001758
16749.000000   1.001937
16999.000000   1.002110
17249.000000   1.001937
17499.000000   1.002289
17749.000000   1.002289
17999.000000   1.002289
18249.000000   1.002462
18499.000000   1.002462
18748.000000   1.002462
18999.000000   1.002462
19249.000000   1.002462
19499.000000   1.002642
19749.000000   1.002642
19999.000000   1.002462
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = No
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 25 October 2019  12:02:56
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 5
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 15:32:54
@@Data
New Section: Section 0: 
2.967100E+1   1.300147E+2   1.300147E+2   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -1.917457E-1   2.789382E-1   -3.002157E-4   -4.054084E-5   4.054084E-5   -3.002157E-4   3.029406E-4   -1.723094E+2   -8.230935E+1   
5.526600E+1   1.299494E+2   1.299494E+2   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -1.760441E-1   2.585904E-1   -2.772559E-4   -3.885142E-5   3.885142E-5   -2.772559E-4   2.799648E-4   -1.720232E+2   -8.202318E+1   
8.030500E+1   1.299950E+2   1.299950E+2   8.998000E+3   8.998000E+3   9.000000E+1   8.998000E+3   8.998000E+3   -1.568365E-1   2.356433E-1   -2.504356E-4   -3.805579E-5   3.805579E-5   -2.504356E-4   2.533106E-4   -1.713595E+2   -8.135953E+1   
1.051670E+2   1.300454E+2   1.300454E+2   8.497000E+3   8.497000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -1.447283E-1   2.171790E-1   -2.309241E-4   -3.493996E-5   3.493996E-5   -2.309241E-4   2.335525E-4   -1.713961E+2   -8.139613E+1   
1.305260E+2   1.300142E+2   1.300142E+2   7.998000E+3   7.998000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -1.279952E-1   1.943023E-1   -2.056797E-4   -3.236017E-5   3.236017E-5   -2.056797E-4   2.082098E-4   -1.710588E+2   -8.105878E+1   
1.563780E+2   1.300107E+2   1.300107E+2   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -1.103381E-1   1.728249E-1   -1.807752E-4   -3.137862E-5   3.137862E-5   -1.807752E-4   1.834783E-4   -1.701528E+2   -8.015282E+1   
1.817150E+2   1.300697E+2   1.300697E+2   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -9.364130E-2   1.506767E-1   -1.560276E-4   -2.924814E-5   2.924814E-5   -1.560276E-4   1.587452E-4   -1.693828E+2   -7.938284E+1   
2.071360E+2   1.300410E+2   1.300410E+2   6.497000E+3   6.497000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -7.898657E-2   1.299982E-1   -1.334997E-4   -2.656826E-5   2.656826E-5   -1.334997E-4   1.361177E-4   -1.687444E+2   -7.874442E+1   
2.326170E+2   1.300559E+2   1.300559E+2   5.998000E+3   5.998000E+3   9.000000E+1   5.998000E+3   5.998000E+3   -5.885207E-2   1.072717E-1   -1.062500E-4   -2.660236E-5   2.660236E-5   -1.062500E-4   1.095297E-4   -1.659435E+2   -7.594353E+1   
2.581970E+2   1.299715E+2   1.299715E+2   5.498000E+3   5.498000E+3   9.000000E+1   5.498000E+3   5.498000E+3   -4.804645E-2   8.948410E-2   -8.798461E-5   -2.296553E-5   2.296553E-5   -8.798461E-5   9.093243E-5   -1.653712E+2   -7.537118E+1   
2.836380E+2   1.300242E+2   1.300242E+2   4.997000E+3   4.997000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -2.980936E-2   6.576655E-2   -6.126260E-5   -2.094839E-5   2.094839E-5   -6.126260E-5   6.474520E-5   -1.611222E+2   -7.112217E+1   
3.088170E+2   1.300449E+2   1.300449E+2   4.498000E+3   4.498000E+3   9.000000E+1   4.498000E+3   4.498000E+3   -1.687153E-2   4.760406E-2   -4.143479E-5   -1.864348E-5   1.864348E-5   -4.143479E-5   4.543590E-5   -1.557747E+2   -6.577475E+1   
3.346730E+2   1.299859E+2   1.299859E+2   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -1.107528E-3   2.764035E-2   -1.868659E-5   -1.725132E-5   1.725132E-5   -1.868659E-5   2.543220E-5   -1.372870E+2   -4.728704E+1   
3.604220E+2   1.300260E+2   1.300260E+2   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   1.104644E-2   7.481481E-3   1.956815E-6   -1.306147E-5   1.306147E-5   1.956815E-6   1.320724E-5   -8.147955E+1   8.520445E+0   
3.858800E+2   1.300769E+2   1.300769E+2   2.998000E+3   2.998000E+3   9.000000E+1   2.998000E+3   2.998000E+3   2.548848E-2   -9.921417E-3   2.221989E-5   -1.236573E-5   1.236573E-5   2.221989E-5   2.542901E-5   -2.909665E+1   6.090335E+1   
4.117310E+2   1.301405E+2   1.301405E+2   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   4.006514E-2   -3.031895E-2   4.451655E-5   -9.811752E-6   9.811752E-6   4.451655E-5   4.558502E-5   -1.242965E+1   7.757035E+1   
4.374800E+2   1.300243E+2   1.300243E+2   1.999000E+3   1.999000E+3   9.000000E+1   1.999000E+3   1.999000E+3   5.383600E-2   -5.105922E-2   6.653826E-5   -6.437707E-6   6.437707E-6   6.653826E-5   6.684897E-5   -5.526278E+0   8.447372E+1   
4.713780E+2   1.300142E+2   1.300142E+2   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   5.540586E-2   -5.180627E-2   6.799537E-5   -7.110418E-6   7.110418E-6   6.799537E-5   6.836614E-5   -5.969842E+0   8.403016E+1   
4.934530E+2   1.300017E+2   1.300017E+2   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   5.690393E-2   -5.386607E-2   7.026307E-5   -6.871796E-6   6.871796E-6   7.026307E-5   7.059831E-5   -5.585818E+0   8.441418E+1   
5.154770E+2   1.299997E+2   1.299997E+2   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   5.800286E-2   -5.477603E-2   7.153513E-5   -7.089697E-6   7.089697E-6   7.153513E-5   7.188559E-5   -5.659981E+0   8.434002E+1   
5.375940E+2   1.300393E+2   1.300393E+2   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   6.136593E-2   -5.836028E-2   7.594872E-5   -7.233847E-6   7.233847E-6   7.594872E-5   7.629244E-5   -5.440807E+0   8.455919E+1   
5.596860E+2   1.299557E+2   1.299557E+2   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   6.121097E-2   -5.934415E-2   7.649370E-5   -6.476009E-6   6.476009E-6   7.649370E-5   7.676735E-5   -4.839160E+0   8.516084E+1   
5.817550E+2   1.300486E+2   1.300486E+2   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   6.256702E-2   -6.094164E-2   7.837250E-5   -6.434588E-6   6.434588E-6   7.837250E-5   7.863621E-5   -4.693606E+0   8.530639E+1   
6.040380E+2   1.299951E+2   1.299951E+2   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   6.492901E-2   -6.290419E-2   8.111098E-5   -6.898534E-6   6.898534E-6   8.111098E-5   8.140381E-5   -4.861339E+0   8.513866E+1   
6.260640E+2   1.299998E+2   1.299998E+2   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   6.650499E-2   -6.531895E-2   8.365804E-5   -6.485472E-6   6.485472E-6   8.365804E-5   8.390905E-5   -4.432909E+0   8.556709E+1   
6.480600E+2   1.300744E+2   1.300744E+2   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   6.695721E-2   -6.699434E-2   8.502879E-5   -5.724625E-6   5.724625E-6   8.502879E-5   8.522128E-5   -3.851667E+0   8.614833E+1   
6.702400E+2   1.299645E+2   1.299645E+2   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   6.837460E-2   -6.986038E-2   8.777170E-5   -4.899230E-6   4.899230E-6   8.777170E-5   8.790833E-5   -3.194813E+0   8.680519E+1   
6.925350E+2   1.300175E+2   1.300175E+2   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   6.941554E-2   -6.987544E-2   8.842506E-5   -5.659305E-6   5.659305E-6   8.842506E-5   8.860598E-5   -3.662001E+0   8.633800E+1   
7.148280E+2   1.300240E+2   1.300240E+2   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   7.094519E-2   -7.361400E-2   9.180566E-5   -4.346513E-6   4.346513E-6   9.180566E-5   9.190849E-5   -2.710629E+0   8.728937E+1   
7.371090E+2   1.300565E+2   1.300565E+2   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   7.162658E-2   -7.450954E-2   9.281018E-5   -4.265016E-6   4.265016E-6   9.281018E-5   9.290812E-5   -2.631130E+0   8.736887E+1   
7.593550E+2   1.299795E+2   1.299795E+2   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   7.303539E-2   -7.671476E-2   9.511741E-5   -3.865306E-6   3.865306E-6   9.511741E-5   9.519591E-5   -2.327060E+0   8.767294E+1   
7.816640E+2   1.299905E+2   1.299905E+2   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   7.430950E-2   -7.828493E-2   9.692776E-5   -3.781140E-6   3.781140E-6   9.692776E-5   9.700148E-5   -2.233969E+0   8.776603E+1   
8.038820E+2   1.300077E+2   1.300077E+2   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   7.601436E-2   -7.910282E-2   9.851446E-5   -4.507396E-6   4.507396E-6   9.851446E-5   9.861752E-5   -2.619664E+0   8.738034E+1   
8.261990E+2   1.300164E+2   1.300164E+2   1.148000E+3   1.148000E+3   9.000000E+1   1.148000E+3   1.148000E+3   7.638833E-2   -8.117368E-2   1.000944E-4   -3.430122E-6   3.430122E-6   1.000944E-4   1.001531E-4   -1.962694E+0   8.803731E+1   
8.484280E+2   1.300772E+2   1.300772E+2   1.097000E+3   1.097000E+3   9.000000E+1   1.098000E+3   1.098000E+3   7.792873E-2   -8.325311E-2   1.024011E-4   -3.209976E-6   3.209976E-6   1.024011E-4   1.024514E-4   -1.795468E+0   8.820453E+1   
8.707050E+2   1.300155E+2   1.300155E+2   1.047000E+3   1.047000E+3   9.000000E+1   1.048000E+3   1.048000E+3   7.923904E-2   -8.396948E-2   1.036777E-4   -3.710786E-6   3.710786E-6   1.036777E-4   1.037441E-4   -2.049830E+0   8.795017E+1   
8.928430E+2   1.299879E+2   1.299879E+2   9.970000E+2   9.970000E+2   9.000000E+1   9.980000E+2   9.980000E+2   7.973298E-2   -8.513193E-2   1.047402E-4   -3.316138E-6   3.316138E-6   1.047402E-4   1.047927E-4   -1.813413E+0   8.818659E+1   
9.147250E+2   1.300384E+2   1.300384E+2   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   8.207473E-2   -8.705950E-2   1.074434E-4   -3.787977E-6   3.787977E-6   1.074434E-4   1.075101E-4   -2.019159E+0   8.798084E+1   
9.366480E+2   1.299441E+2   1.299441E+2   8.970000E+2   8.970000E+2   9.000000E+1   8.980000E+2   8.980000E+2   8.228857E-2   -8.906101E-2   1.088791E-4   -2.637610E-6   2.637610E-6   1.088791E-4   1.089111E-4   -1.387726E+0   8.861227E+1   
9.585350E+2   1.300586E+2   1.300586E+2   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   8.347186E-2   -9.127701E-2   1.110540E-4   -2.064050E-6   2.064050E-6   1.110540E-4   1.110731E-4   -1.064777E+0   8.893522E+1   
9.803610E+2   1.300319E+2   1.300319E+2   7.970000E+2   7.970000E+2   9.000000E+1   7.980000E+2   7.980000E+2   8.462294E-2   -9.342865E-2   1.131669E-4   -1.508740E-6   1.508740E-6   1.131669E-4   1.131770E-4   -7.638210E-1   8.923618E+1   
1.002287E+3   1.300258E+2   1.300258E+2   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   8.539114E-2   -9.439512E-2   1.142713E-4   -1.445081E-6   1.445081E-6   1.142713E-4   1.142805E-4   -7.245268E-1   8.927547E+1   
1.024183E+3   1.300015E+2   1.300015E+2   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   8.714387E-2   -9.665632E-2   1.168277E-4   -1.263144E-6   1.263144E-6   1.168277E-4   1.168345E-4   -6.194594E-1   8.938054E+1   
1.046006E+3   1.300036E+2   1.300036E+2   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   8.768871E-2   -9.824919E-2   1.182019E-4   -6.247507E-7   6.247507E-7   1.182019E-4   1.182036E-4   -3.028313E-1   8.969717E+1   
1.067881E+3   1.300349E+2   1.300349E+2   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   8.976945E-2   -1.004354E-1   1.209122E-4   -7.344313E-7   7.344313E-7   1.209122E-4   1.209144E-4   -3.480153E-1   8.965198E+1   
1.089757E+3   1.300178E+2   1.300178E+2   5.480000E+2   5.480000E+2   9.000000E+1   5.480000E+2   5.480000E+2   9.077758E-2   -1.014107E-1   1.221707E-4   -8.424715E-7   8.424715E-7   1.221707E-4   1.221736E-4   -3.950973E-1   8.960490E+1   
1.111594E+3   1.300119E+2   1.300119E+2   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   9.160038E-2   -1.039273E-1   1.243184E-4   1.942539E-7   -1.942539E-7   1.243184E-4   1.243185E-4   8.952754E-2   9.008953E+1   
1.133468E+3   1.300509E+2   1.300509E+2   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   9.202134E-2   -1.065611E-1   1.262940E-4   1.604821E-6   -1.604821E-6   1.262940E-4   1.263042E-4   7.280196E-1   9.072802E+1   
1.155240E+3   1.300309E+2   1.300309E+2   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   9.310678E-2   -1.071057E-1   1.273198E-4   1.158011E-6   -1.158011E-6   1.273198E-4   1.273250E-4   5.211079E-1   9.052111E+1   
1.177116E+3   1.300083E+2   1.300083E+2   3.480000E+2   3.480000E+2   9.000000E+1   3.480000E+2   3.480000E+2   9.537751E-2   -1.091851E-1   1.300779E-4   8.379735E-7   -8.379735E-7   1.300779E-4   1.300806E-4   3.690993E-1   9.036910E+1   
1.199002E+3   1.301138E+2   1.301138E+2   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   9.714071E-2   -1.105098E-1   1.320308E-4   3.999253E-7   -3.999253E-7   1.320308E-4   1.320314E-4   1.735501E-1   9.017355E+1   
1.220879E+3   1.300880E+2   1.300880E+2   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   9.821081E-2   -1.121374E-1   1.337524E-4   6.724906E-7   -6.724906E-7   1.337524E-4   1.337541E-4   2.880737E-1   9.028807E+1   
1.242663E+3   1.300050E+2   1.300050E+2   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   9.880755E-2   -1.144472E-1   1.356257E-4   1.741218E-6   -1.741218E-6   1.356257E-4   1.356369E-4   7.355459E-1   9.073555E+1   
1.264547E+3   1.300083E+2   1.300083E+2   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   1.002231E-1   -1.154348E-1   1.371441E-4   1.339887E-6   -1.339887E-6   1.371441E-4   1.371506E-4   5.597576E-1   9.055976E+1   
1.286422E+3   1.300346E+2   1.300346E+2   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   1.014076E-1   -1.168147E-1   1.387751E-4   1.365965E-6   -1.365965E-6   1.387751E-4   1.387818E-4   5.639449E-1   9.056394E+1   
1.308168E+3   1.299155E+2   1.299155E+2   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   1.025860E-1   -1.197998E-1   1.414478E-4   2.445948E-6   -2.445948E-6   1.414478E-4   1.414690E-4   9.906728E-1   9.099067E+1   
1.341343E+3   1.299868E+2   1.299868E+2   4.700000E+1   4.700000E+1   9.000000E+1   4.700000E+1   4.700000E+1   1.036766E-1   -1.182984E-1   1.411442E-4   6.576851E-7   -6.576851E-7   1.411442E-4   1.411458E-4   2.669773E-1   9.026698E+1   
1.362777E+3   1.300107E+2   1.300107E+2   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   1.017328E-1   -1.193642E-1   1.406366E-4   2.792181E-6   -2.792181E-6   1.406366E-4   1.406643E-4   1.137393E+0   9.113739E+1   
1.381842E+3   1.300646E+2   1.300646E+2   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   1.042786E-1   -1.180612E-1   1.413619E-4   5.742641E-8   -5.742641E-8   1.413619E-4   1.413619E-4   2.327565E-2   9.002328E+1   
1.404273E+3   1.300834E+2   1.300834E+2   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   1.019586E-1   -1.201404E-1   1.412817E-4   3.132636E-6   -3.132636E-6   1.412817E-4   1.413165E-4   1.270209E+0   9.127021E+1   
1.423356E+3   1.299971E+2   1.299971E+2   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   1.023648E-1   -1.197606E-1   1.412855E-4   2.583881E-6   -2.583881E-6   1.412855E-4   1.413091E-4   1.047729E+0   9.104773E+1   
1.445787E+3   1.300104E+2   1.300104E+2   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   1.038402E-1   -1.189049E-1   1.416404E-4   9.332619E-7   -9.332619E-7   1.416404E-4   1.416434E-4   3.775138E-1   9.037751E+1   
1.464917E+3   1.300994E+2   1.300994E+2   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   1.034116E-1   -1.196523E-1   1.418621E-4   1.738848E-6   -1.738848E-6   1.418621E-4   1.418728E-4   7.022571E-1   9.070226E+1   
1.487327E+3   1.299651E+2   1.299651E+2   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   1.027808E-1   -1.210331E-1   1.423715E-4   3.108155E-6   -3.108155E-6   1.423715E-4   1.424054E-4   1.250642E+0   9.125064E+1   
1.506338E+3   1.300092E+2   1.300092E+2   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   1.038150E-1   -1.199278E-1   1.422910E-4   1.620580E-6   -1.620580E-6   1.422910E-4   1.423002E-4   6.525245E-1   9.065252E+1   
1.528833E+3   1.300555E+2   1.300555E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   1.035757E-1   -1.192743E-1   1.417174E-4   1.370334E-6   -1.370334E-6   1.417174E-4   1.417241E-4   5.540033E-1   9.055400E+1   
1.547850E+3   1.299535E+2   1.299535E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   1.030799E-1   -1.197995E-1   1.417530E-4   2.080417E-6   -2.080417E-6   1.417530E-4   1.417683E-4   8.408325E-1   9.084083E+1   
1.570239E+3   1.299816E+2   1.299816E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   1.036310E-1   -1.192004E-1   1.417034E-4   1.281166E-6   -1.281166E-6   1.417034E-4   1.417092E-4   5.180072E-1   9.051801E+1   
1.589277E+3   1.300152E+2   1.300152E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   1.041215E-1   -1.186303E-1   1.416355E-4   5.456704E-7   -5.456704E-7   1.416355E-4   1.416365E-4   2.207389E-1   9.022074E+1   
1.611695E+3   1.300144E+2   1.300144E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   1.035429E-1   -1.209742E-1   1.428043E-4   2.505994E-6   -2.505994E-6   1.428043E-4   1.428263E-4   1.005349E+0   9.100535E+1   
1.630708E+3   1.300442E+2   1.300442E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   1.029296E-1   -1.207331E-1   1.422681E-4   2.801942E-6   -2.801942E-6   1.422681E-4   1.422957E-4   1.128283E+0   9.112828E+1   
1.653097E+3   1.300571E+2   1.300571E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   1.039500E-1   -1.199486E-1   1.423880E-4   1.534373E-6   -1.534373E-6   1.423880E-4   1.423963E-4   6.173952E-1   9.061740E+1   
1.672158E+3   1.300556E+2   1.300556E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   1.019718E-1   -1.206941E-1   1.416506E-4   3.484905E-6   -3.484905E-6   1.416506E-4   1.416934E-4   1.409314E+0   9.140931E+1   
1.694580E+3   1.300011E+2   1.300011E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   1.031984E-1   -1.205702E-1   1.423281E-4   2.496665E-6   -2.496665E-6   1.423281E-4   1.423500E-4   1.004957E+0   9.100496E+1   
1.713591E+3   1.299752E+2   1.299752E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   1.045633E-1   -1.196645E-1   1.425822E-4   8.950359E-7   -8.950359E-7   1.425822E-4   1.425850E-4   3.596600E-1   9.035966E+1   
1.735669E+3   1.299794E+2   1.299794E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   1.045709E-1   -1.206125E-1   1.432043E-4   1.509143E-6   -1.509143E-6   1.432043E-4   1.432123E-4   6.037830E-1   9.060378E+1   
1.754421E+3   1.300383E+2   1.300383E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   1.028750E-1   -1.207040E-1   1.422154E-4   2.823294E-6   -2.823294E-6   1.422154E-4   1.422434E-4   1.137301E+0   9.113730E+1   
1.776433E+3   1.300678E+2   1.300678E+2   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   1.047023E-1   -1.211675E-1   1.436470E-4   1.774866E-6   -1.774866E-6   1.436470E-4   1.436579E-4   7.078964E-1   9.070790E+1   
1.795141E+3   1.299779E+2   1.299779E+2   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   1.030625E-1   -1.206693E-1   1.423087E-4   2.661967E-6   -2.661967E-6   1.423087E-4   1.423336E-4   1.071626E+0   9.107163E+1   
1.817175E+3   1.300068E+2   1.300068E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   1.045038E-1   -1.208368E-1   1.433088E-4   1.705444E-6   -1.705444E-6   1.433088E-4   1.433190E-4   6.818151E-1   9.068182E+1   
1.835896E+3   1.300059E+2   1.300059E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   1.039000E-1   -1.207469E-1   1.428770E-4   2.093251E-6   -2.093251E-6   1.428770E-4   1.428924E-4   8.393644E-1   9.083936E+1   
1.857976E+3   1.299699E+2   1.299699E+2   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   1.048900E-1   -1.211083E-1   1.437245E-4   1.597281E-6   -1.597281E-6   1.437245E-4   1.437334E-4   6.367299E-1   9.063673E+1   
1.880001E+3   1.300409E+2   1.300409E+2   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   1.046056E-1   -1.227895E-1   1.446436E-4   2.906741E-6   -2.906741E-6   1.446436E-4   1.446728E-4   1.151254E+0   9.115125E+1   
1.902086E+3   1.300266E+2   1.300266E+2   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   1.045314E-1   -1.212221E-1   1.435769E-4   1.936954E-6   -1.936954E-6   1.435769E-4   1.435899E-4   7.729137E-1   9.077291E+1   
1.924104E+3   1.300120E+2   1.300120E+2   -8.000000E+0   -8.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   1.045209E-1   -1.216627E-1   1.438574E-4   2.232685E-6   -2.232685E-6   1.438574E-4   1.438747E-4   8.891667E-1   9.088917E+1   
1.946175E+3   1.300344E+2   1.300344E+2   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   1.045489E-1   -1.224011E-1   1.443555E-4   2.694798E-6   -2.694798E-6   1.443555E-4   1.443807E-4   1.069461E+0   9.106946E+1   
1.968386E+3   1.300096E+2   1.300096E+2   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   1.053162E-1   -1.219219E-1   1.445178E-4   1.814007E-6   -1.814007E-6   1.445178E-4   1.445292E-4   7.191465E-1   9.071915E+1   
1.990660E+3   1.299914E+2   1.299914E+2   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   1.038868E-1   -1.214292E-1   1.433132E-4   2.549068E-6   -2.549068E-6   1.433132E-4   1.433359E-4   1.018995E+0   9.101899E+1   
2.012933E+3   1.300204E+2   1.300204E+2   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   1.056708E-1   -1.218633E-1   1.446989E-4   1.513380E-6   -1.513380E-6   1.446989E-4   1.447068E-4   5.992246E-1   9.059922E+1   
2.035204E+3   1.299727E+2   1.299727E+2   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   1.049011E-1   -1.212200E-1   1.438040E-4   1.662115E-6   -1.662115E-6   1.438040E-4   1.438137E-4   6.622061E-1   9.066221E+1   
2.057490E+3   1.300064E+2   1.300064E+2   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   1.050437E-1   -1.219698E-1   1.443806E-4   2.046804E-6   -2.046804E-6   1.443806E-4   1.443951E-4   8.121964E-1   9.081220E+1   
2.079760E+3   1.300713E+2   1.300713E+2   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   1.051376E-1   -1.230709E-1   1.451557E-4   2.697218E-6   -2.697218E-6   1.451557E-4   1.451808E-4   1.064522E+0   9.106452E+1   
2.101996E+3   1.299964E+2   1.299964E+2   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   1.061967E-1   -1.212602E-1   1.446312E-4   7.301193E-7   -7.301193E-7   1.446312E-4   1.446331E-4   2.892349E-1   9.028923E+1   
2.124233E+3   1.300166E+2   1.300166E+2   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   1.043390E-1   -1.228858E-1   1.445415E-4   3.166915E-6   -3.166915E-6   1.445415E-4   1.445762E-4   1.255154E+0   9.125515E+1   
2.146469E+3   1.299598E+2   1.299598E+2   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   1.049713E-1   -1.226162E-1   1.447568E-4   2.522955E-6   -2.522955E-6   1.447568E-4   1.447788E-4   9.985027E-1   9.099850E+1   
2.168740E+3   1.300072E+2   1.300072E+2   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   1.042872E-1   -1.224898E-1   1.442515E-4   2.946336E-6   -2.946336E-6   1.442515E-4   1.442816E-4   1.170103E+0   9.117010E+1   
2.191016E+3   1.300243E+2   1.300243E+2   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   1.056205E-1   -1.214252E-1   1.443825E-4   1.264186E-6   -1.264186E-6   1.443825E-4   1.443880E-4   5.016583E-1   9.050166E+1   
2.213245E+3   1.299757E+2   1.299757E+2   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   1.049477E-1   -1.227763E-1   1.448465E-4   2.645120E-6   -2.645120E-6   1.448465E-4   1.448706E-4   1.046193E+0   9.104619E+1   
2.235477E+3   1.299791E+2   1.299791E+2   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   1.044820E-1   -1.233985E-1   1.449638E-4   3.396342E-6   -3.396342E-6   1.449638E-4   1.450036E-4   1.342132E+0   9.134213E+1   
2.257753E+3   1.299689E+2   1.299689E+2   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   1.060657E-1   -1.225515E-1   1.453912E-4   1.671220E-6   -1.671220E-6   1.453912E-4   1.454008E-4   6.585656E-1   9.065857E+1   
2.280002E+3   1.300778E+2   1.300778E+2   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   1.057248E-1   -1.225223E-1   1.451615E-4   1.904275E-6   -1.904275E-6   1.451615E-4   1.451740E-4   7.515814E-1   9.075158E+1   
2.302271E+3   1.300154E+2   1.300154E+2   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   1.036343E-1   -1.229248E-1   1.441312E-4   3.713623E-6   -3.713623E-6   1.441312E-4   1.441790E-4   1.475932E+0   9.147593E+1   
2.324550E+3   1.300390E+2   1.300390E+2   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   1.063730E-1   -1.235556E-1   1.462352E-4   2.100342E-6   -2.100342E-6   1.462352E-4   1.462503E-4   8.228692E-1   9.082287E+1   
2.346839E+3   1.299881E+2   1.299881E+2   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   1.067458E-1   -1.238495E-1   1.466571E-4   2.016793E-6   -2.016793E-6   1.466571E-4   1.466710E-4   7.878682E-1   9.078787E+1   
2.369087E+3   1.300346E+2   1.300346E+2   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   1.057969E-1   -1.225389E-1   1.452169E-4   1.861786E-6   -1.861786E-6   1.452169E-4   1.452288E-4   7.345336E-1   9.073453E+1   
2.391356E+3   1.299848E+2   1.299848E+2   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   1.050449E-1   -1.230417E-1   1.450795E-4   2.746689E-6   -2.746689E-6   1.450795E-4   1.451055E-4   1.084612E+0   9.108461E+1   
2.424692E+3   1.300254E+2   1.300254E+2   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   1.083703E-1   -1.251113E-1   1.484833E-4   1.640229E-6   -1.640229E-6   1.484833E-4   1.484923E-4   6.328953E-1   9.063290E+1   
2.446373E+3   1.300329E+2   1.300329E+2   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   1.082433E-1   -1.261992E-1   1.491133E-4   2.445409E-6   -2.445409E-6   1.491133E-4   1.491333E-4   9.395480E-1   9.093955E+1   
2.468103E+3   1.300382E+2   1.300382E+2   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   1.094416E-1   -1.287882E-1   1.515403E-4   3.251721E-6   -3.251721E-6   1.515403E-4   1.515752E-4   1.229252E+0   9.122925E+1   
2.489882E+3   1.300792E+2   1.300792E+2   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   1.110440E-1   -1.302440E-1   1.534791E-4   3.018250E-6   -3.018250E-6   1.534791E-4   1.535088E-4   1.126608E+0   9.112661E+1   
2.511570E+3   1.300459E+2   1.300459E+2   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   1.109341E-1   -1.311702E-1   1.540144E-4   3.705023E-6   -3.705023E-6   1.540144E-4   1.540590E-4   1.378061E+0   9.137806E+1   
2.533350E+3   1.300727E+2   1.300727E+2   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   1.115839E-1   -1.325151E-1   1.552921E-4   4.103729E-6   -4.103729E-6   1.552921E-4   1.553463E-4   1.513739E+0   9.151374E+1   
2.555035E+3   1.300054E+2   1.300054E+2   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   1.139490E-1   -1.342047E-1   1.578547E-4   3.458999E-6   -3.458999E-6   1.578547E-4   1.578926E-4   1.255296E+0   9.125530E+1   
2.576731E+3   1.299835E+2   1.299835E+2   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   1.148056E-1   -1.361912E-1   1.596780E-4   4.124166E-6   -4.124166E-6   1.596780E-4   1.597313E-4   1.479507E+0   9.147951E+1   
2.598470E+3   1.300608E+2   1.300608E+2   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   1.154658E-1   -1.373376E-1   1.608329E-4   4.385375E-6   -4.385375E-6   1.608329E-4   1.608927E-4   1.561877E+0   9.156188E+1   
2.620109E+3   1.300623E+2   1.300623E+2   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   1.171639E-1   -1.396447E-1   1.633853E-4   4.637730E-6   -4.637730E-6   1.633853E-4   1.634511E-4   1.625917E+0   9.162592E+1   
2.641845E+3   1.300435E+2   1.300435E+2   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   1.167623E-1   -1.402770E-1   1.635488E-4   5.348139E-6   -5.348139E-6   1.635488E-4   1.636363E-4   1.872937E+0   9.187294E+1   
2.663482E+3   1.299512E+2   1.299512E+2   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.490000E+2   -6.490000E+2   1.182720E-1   -1.422448E-1   1.657638E-4   5.517973E-6   -5.517973E-6   1.657638E-4   1.658556E-4   1.906568E+0   9.190657E+1   
2.685186E+3   1.300119E+2   1.300119E+2   -7.010000E+2   -7.010000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   1.190605E-1   -1.432949E-1   1.669352E-4   5.621365E-6   -5.621365E-6   1.669352E-4   1.670298E-4   1.928645E+0   9.192865E+1   
2.706845E+3   1.300317E+2   1.300317E+2   -7.500000E+2   -7.500000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   1.208672E-1   -1.454544E-1   1.694587E-4   5.696894E-6   -5.696894E-6   1.694587E-4   1.695544E-4   1.925455E+0   9.192546E+1   
2.728533E+3   1.300153E+2   1.300153E+2   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   1.214817E-1   -1.461325E-1   1.702802E-4   5.685659E-6   -5.685659E-6   1.702802E-4   1.703751E-4   1.912397E+0   9.191240E+1   
2.750160E+3   1.300389E+2   1.300389E+2   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   1.234028E-1   -1.478054E-1   1.725575E-4   5.358435E-6   -5.358435E-6   1.725575E-4   1.726407E-4   1.778637E+0   9.177864E+1   
2.771877E+3   1.300095E+2   1.300095E+2   -9.000000E+2   -9.000000E+2   9.000000E+1   -9.000000E+2   -9.000000E+2   1.228030E-1   -1.495483E-1   1.733218E-4   6.941510E-6   -6.941510E-6   1.733218E-4   1.734607E-4   2.293461E+0   9.229346E+1   
2.793584E+3   1.299892E+2   1.299892E+2   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   1.245646E-1   -1.513255E-1   1.755684E-4   6.800501E-6   -6.800501E-6   1.755684E-4   1.757000E-4   2.218197E+0   9.221820E+1   
2.815269E+3   1.300158E+2   1.300158E+2   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   1.255271E-1   -1.526500E-1   1.770260E-4   6.954529E-6   -6.954529E-6   1.770260E-4   1.771626E-4   2.249728E+0   9.224973E+1   
2.837354E+3   1.299973E+2   1.299973E+2   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   1.265563E-1   -1.537112E-1   1.783535E-4   6.887027E-6   -6.887027E-6   1.783535E-4   1.784864E-4   2.211348E+0   9.221135E+1   
2.859223E+3   1.299652E+2   1.299652E+2   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   1.277292E-1   -1.550791E-1   1.799696E-4   6.913869E-6   -6.913869E-6   1.799696E-4   1.801023E-4   2.200043E+0   9.220004E+1   
2.881098E+3   1.299914E+2   1.299914E+2   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   1.285870E-1   -1.571500E-1   1.818486E-4   7.633297E-6   -7.633297E-6   1.818486E-4   1.820087E-4   2.403643E+0   9.240364E+1   
2.903667E+3   1.300102E+2   1.300102E+2   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   1.297586E-1   -1.586410E-1   1.835441E-4   7.741486E-6   -7.741486E-6   1.835441E-4   1.837073E-4   2.415179E+0   9.241518E+1   
2.925446E+3   1.300317E+2   1.300317E+2   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.250000E+3   -1.250000E+3   1.300473E-1   -1.615166E-1   1.855954E-4   9.407929E-6   -9.407929E-6   1.855954E-4   1.858337E-4   2.901870E+0   9.290187E+1   
2.947327E+3   1.300136E+2   1.300136E+2   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   1.320721E-1   -1.616884E-1   1.869591E-4   8.022627E-6   -8.022627E-6   1.869591E-4   1.871312E-4   2.457120E+0   9.245712E+1   
2.969930E+3   1.299719E+2   1.299719E+2   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   1.323550E-1   -1.638157E-1   1.885195E-4   9.204167E-6   -9.204167E-6   1.885195E-4   1.887440E-4   2.795157E+0   9.279516E+1   
2.991731E+3   1.300337E+2   1.300337E+2   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   1.355797E-1   -1.653343E-1   1.915022E-4   7.811927E-6   -7.811927E-6   1.915022E-4   1.916615E-4   2.335965E+0   9.233596E+1   
3.013858E+3   1.299740E+2   1.299740E+2   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   1.358417E-1   -1.683037E-1   1.935981E-4   9.559489E-6   -9.559489E-6   1.935981E-4   1.938340E-4   2.826855E+0   9.282686E+1   
3.036177E+3   1.300231E+2   1.300231E+2   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   1.369680E-1   -1.691858E-1   1.948689E-4   9.303138E-6   -9.303138E-6   1.948689E-4   1.950908E-4   2.733254E+0   9.273325E+1   
3.058277E+3   1.300374E+2   1.300374E+2   -1.550000E+3   -1.550000E+3   9.000000E+1   -1.548000E+3   -1.548000E+3   1.384485E-1   -1.717711E-1   1.974681E-4   9.898259E-6   -9.898259E-6   1.974681E-4   1.977160E-4   2.869599E+0   9.286960E+1   
3.080315E+3   1.299577E+2   1.299577E+2   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   1.390115E-1   -1.739846E-1   1.992578E-4   1.092902E-5   -1.092902E-5   1.992578E-4   1.995572E-4   3.139451E+0   9.313945E+1   
3.103197E+3   1.300470E+2   1.300470E+2   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   1.419383E-1   -1.768547E-1   2.029365E-4   1.064062E-5   -1.064062E-5   2.029365E-4   2.032152E-4   3.001455E+0   9.300145E+1   
3.125265E+3   1.300662E+2   1.300662E+2   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.698000E+3   -1.698000E+3   1.417055E-1   -1.775180E-1   2.032245E-4   1.124648E-5   -1.124648E-5   2.032245E-4   2.035355E-4   3.167527E+0   9.316753E+1   
3.147330E+3   1.300072E+2   1.300072E+2   -1.750000E+3   -1.750000E+3   9.000000E+1   -1.748000E+3   -1.748000E+3   1.428078E-1   -1.802199E-1   2.056657E-4   1.219761E-5   -1.219761E-5   2.056657E-4   2.060271E-4   3.394119E+0   9.339412E+1   
3.170473E+3   1.300402E+2   1.300402E+2   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.798000E+3   -1.798000E+3   1.463015E-1   -1.806175E-1   2.080847E-4   9.873473E-6   -9.873473E-6   2.080847E-4   2.083188E-4   2.716607E+0   9.271661E+1   
3.192530E+3   1.300289E+2   1.300289E+2   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.848000E+3   -1.848000E+3   1.454253E-1   -1.831203E-1   2.091730E-4   1.215780E-5   -1.215780E-5   2.091730E-4   2.095260E-4   3.326471E+0   9.332647E+1   
3.214650E+3   1.300227E+2   1.300227E+2   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   1.487460E-1   -1.849942E-1   2.124465E-4   1.092682E-5   -1.092682E-5   2.124465E-4   2.127274E-4   2.944314E+0   9.294431E+1   
3.237993E+3   1.300631E+2   1.300631E+2   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   1.488356E-1   -1.870769E-1   2.138583E-4   1.222214E-5   -1.222214E-5   2.138583E-4   2.142073E-4   3.270932E+0   9.327093E+1   
3.259809E+3   1.300435E+2   1.300435E+2   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   1.492648E-1   -1.873518E-1   2.143027E-4   1.208441E-5   -1.208441E-5   2.143027E-4   2.146432E-4   3.227459E+0   9.322746E+1   
3.296878E+3   1.300167E+2   1.300167E+2   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.608803E-1   -2.056175E-1   2.333802E-4   1.543485E-5   -1.543485E-5   2.333802E-4   2.338901E-4   3.783807E+0   9.378381E+1   
3.322541E+3   1.299808E+2   1.299808E+2   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.718355E-1   -2.228454E-1   2.513736E-4   1.859516E-5   -1.859516E-5   2.513736E-4   2.520605E-4   4.230702E+0   9.423070E+1   
3.347684E+3   1.299648E+2   1.299648E+2   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.852605E-1   -2.416077E-1   2.718932E-4   2.093181E-5   -2.093181E-5   2.718932E-4   2.726978E-4   4.402255E+0   9.440226E+1   
3.373374E+3   1.299954E+2   1.299954E+2   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   1.937087E-1   -2.557560E-1   2.863310E-4   2.393308E-5   -2.393308E-5   2.863310E-4   2.873295E-4   4.777982E+0   9.477798E+1   
3.399560E+3   1.300142E+2   1.300142E+2   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   1.964352E-1   -2.636722E-1   2.931723E-4   2.709188E-5   -2.709188E-5   2.931723E-4   2.944214E-4   5.279674E+0   9.527967E+1   
3.424321E+3   1.300252E+2   1.300252E+2   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   1.867839E-1   -2.562273E-1   2.823567E-4   2.936298E-5   -2.936298E-5   2.823567E-4   2.838793E-4   5.936993E+0   9.593699E+1   
3.449516E+3   1.300552E+2   1.300552E+2   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   1.722617E-1   -2.377598E-1   2.613507E-4   2.803059E-5   -2.803059E-5   2.613507E-4   2.628496E-4   6.121731E+0   9.612173E+1   
3.475677E+3   1.300271E+2   1.300271E+2   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   1.574203E-1   -2.222303E-1   2.420608E-4   2.885497E-5   -2.885497E-5   2.420608E-4   2.437746E-4   6.797892E+0   9.679789E+1   
3.500357E+3   1.300392E+2   1.300392E+2   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.442739E-1   -2.110410E-1   2.266456E-4   3.126317E-5   -3.126317E-5   2.266456E-4   2.287917E-4   7.853735E+0   9.785373E+1   
3.525007E+3   1.299802E+2   1.299802E+2   -7.001000E+3   -7.001000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.418024E-1   -2.105464E-1   2.247955E-4   3.276784E-5   -3.276784E-5   2.247955E-4   2.271712E-4   8.293440E+0   9.829344E+1   
3.550202E+3   1.300505E+2   1.300505E+2   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.460683E-1   -2.175683E-1   2.320062E-4   3.420334E-5   -3.420334E-5   2.320062E-4   2.345139E-4   8.386378E+0   9.838638E+1   
3.575388E+3   1.299963E+2   1.299963E+2   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.532878E-1   -2.287760E-1   2.437691E-4   3.619092E-5   -3.619092E-5   2.437691E-4   2.464410E-4   8.444673E+0   9.844467E+1   
3.600583E+3   1.300094E+2   1.300094E+2   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.629591E-1   -2.405765E-1   2.574339E-4   3.675252E-5   -3.675252E-5   2.574339E-4   2.600441E-4   8.124922E+0   9.812492E+1   
3.626289E+3   1.300465E+2   1.300465E+2   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.741015E-1   -2.584906E-1   2.759899E-4   4.022300E-5   -4.022300E-5   2.759899E-4   2.789056E-4   8.291956E+0   9.829196E+1   
3.651923E+3   1.299880E+2   1.299880E+2   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.857292E-1   -2.744538E-1   2.935753E-4   4.205911E-5   -4.205911E-5   2.935753E-4   2.965728E-4   8.153011E+0   9.815301E+1   
3.677088E+3   1.299345E+2   1.299345E+2   -1.000000E+4   -1.000000E+4   9.000000E+1   -9.999000E+3   -9.999000E+3   1.991070E-1   -2.929079E-1   3.138651E-4   4.422915E-5   -4.422915E-5   3.138651E-4   3.169661E-4   8.021175E+0   9.802117E+1   
3.713617E+3   1.299929E+2   1.299929E+2   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.823964E-1   -2.697913E-1   2.884782E-4   4.147590E-5   -4.147590E-5   2.884782E-4   2.914445E-4   8.181624E+0   9.818162E+1   
3.738324E+3   1.300207E+2   1.300207E+2   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.665529E-1   -2.483102E-1   2.646925E-4   3.915049E-5   -3.915049E-5   2.646925E-4   2.675722E-4   8.413577E+0   9.841358E+1   
3.762993E+3   1.299934E+2   1.299934E+2   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.500000E+3   -8.500000E+3   1.538707E-1   -2.320658E-1   2.462720E-4   3.791050E-5   -3.791050E-5   2.462720E-4   2.491729E-4   8.751275E+0   9.875127E+1   
3.787593E+3   1.300449E+2   1.300449E+2   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.999000E+3   -7.999000E+3   1.391523E-1   -2.112573E-1   2.236201E-4   3.519266E-5   -3.519266E-5   2.236201E-4   2.263724E-4   8.943683E+0   9.894368E+1   
3.812336E+3   1.300503E+2   1.300503E+2   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.242950E-1   -1.928719E-1   2.024604E-4   3.416176E-5   -3.416176E-5   2.024604E-4   2.053222E-4   9.577479E+0   9.957748E+1   
3.837484E+3   1.300202E+2   1.300202E+2   -7.000000E+3   -7.000000E+3   9.000000E+1   -6.999000E+3   -6.999000E+3   1.122316E-1   -1.738785E-1   1.826320E-4   3.066688E-5   -3.066688E-5   1.826320E-4   1.851889E-4   9.531969E+0   9.953197E+1   
3.862617E+3   1.300351E+2   1.300351E+2   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.003556E-1   -1.556455E-1   1.634148E-4   2.753050E-5   -2.753050E-5   1.634148E-4   1.657176E-4   9.562830E+0   9.956283E+1   
3.886848E+3   1.300603E+2   1.300603E+2   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   8.560530E-2   -1.354564E-1   1.411465E-4   2.524122E-5   -2.524122E-5   1.411465E-4   1.433857E-4   1.013902E+1   1.001390E+2   
3.911593E+3   1.299987E+2   1.299987E+2   -5.499000E+3   -5.499000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   7.508385E-2   -1.178879E-1   1.231995E-4   2.153744E-5   -2.153744E-5   1.231995E-4   1.250679E-4   9.916105E+0   9.991610E+1   
3.936745E+3   1.299767E+2   1.299767E+2   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   6.301217E-2   -1.008735E-1   1.046549E-4   1.934248E-5   -1.934248E-5   1.046549E-4   1.064274E-4   1.047133E+1   1.004713E+2   
3.961021E+3   1.299521E+2   1.299521E+2   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   5.241462E-2   -8.412471E-2   8.719470E-5   1.623088E-5   -1.623088E-5   8.719470E-5   8.869249E-5   1.054465E+1   1.005447E+2   
3.985717E+3   1.300331E+2   1.300331E+2   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   3.910734E-2   -6.673265E-2   6.764025E-5   1.470291E-5   -1.470291E-5   6.764025E-5   6.921979E-5   1.226357E+1   1.022636E+2   
4.010436E+3   1.300625E+2   1.300625E+2   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   2.907704E-2   -4.883741E-2   4.978407E-5   1.042224E-5   -1.042224E-5   4.978407E-5   5.086331E-5   1.182404E+1   1.018240E+2   
4.035072E+3   1.299888E+2   1.299888E+2   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.680312E-2   -3.091138E-2   3.052073E-5   7.780877E-6   -7.780877E-6   3.052073E-5   3.149694E-5   1.430219E+1   1.043022E+2   
4.060194E+3   1.300716E+2   1.300716E+2   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   5.088487E-3   -1.185453E-2   1.086667E-5   3.986556E-6   -3.986556E-6   1.086667E-5   1.157485E-5   2.014611E+1   1.101461E+2   
4.084892E+3   1.300021E+2   1.300021E+2   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.999000E+3   -1.999000E+3   -8.511393E-3   4.669715E-3   -8.303477E-6   3.242363E-6   -3.242363E-6   -8.303477E-6   8.914071E-6   1.586702E+2   2.486702E+2   
4.118557E+3   1.299684E+2   1.299684E+2   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   -8.782904E-3   7.570761E-3   -1.036076E-5   1.546559E-6   -1.546559E-6   -1.036076E-5   1.047555E-5   1.715101E+2   2.615101E+2   
4.140586E+3   1.300758E+2   1.300758E+2   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.899000E+3   -1.899000E+3   -9.103201E-3   1.048101E-2   -1.245420E-5   -1.191803E-7   1.191803E-7   -1.245420E-5   1.245477E-5   -1.794517E+2   -8.945173E+1   
4.162720E+3   1.299770E+2   1.299770E+2   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.849000E+3   -1.849000E+3   -1.160971E-2   1.170543E-2   -1.480129E-5   9.342252E-7   -9.342252E-7   -1.480129E-5   1.483075E-5   1.763884E+2   2.663884E+2   
4.184595E+3   1.299984E+2   1.299984E+2   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.799000E+3   -1.799000E+3   -1.123481E-2   1.262857E-2   -1.517074E-5   5.340833E-8   -5.340833E-8   -1.517074E-5   1.517083E-5   1.797983E+2   2.697983E+2   
4.206673E+3   1.300024E+2   1.300024E+2   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   -1.278504E-2   1.678379E-2   -1.883541E-5   -1.516555E-6   1.516555E-6   -1.883541E-5   1.889637E-5   -1.753967E+2   -8.539669E+1   
4.228709E+3   1.300260E+2   1.300260E+2   -1.700000E+3   -1.700000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   -1.436350E-2   1.679851E-2   -1.982088E-5   -3.587048E-7   3.587048E-7   -1.982088E-5   1.982413E-5   -1.789632E+2   -8.896321E+1   
4.250479E+3   1.301051E+2   1.301051E+2   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   -1.548636E-2   1.965077E-2   -2.237273E-5   -1.392927E-6   1.392927E-6   -2.237273E-5   2.241605E-5   -1.764374E+2   -8.643736E+1   
4.272344E+3   1.301060E+2   1.301060E+2   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.599000E+3   -1.599000E+3   -1.622420E-2   1.982135E-2   -2.293999E-5   -9.587176E-7   9.587176E-7   -2.293999E-5   2.296002E-5   -1.776069E+2   -8.760686E+1   
4.294427E+3   1.300689E+2   1.300689E+2   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   -1.765140E-2   2.253956E-2   -2.559270E-5   -1.680201E-6   1.680201E-6   -2.559270E-5   2.564779E-5   -1.762438E+2   -8.624383E+1   
4.316474E+3   1.300824E+2   1.300824E+2   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   -1.835304E-2   2.489729E-2   -2.756204E-5   -2.702667E-6   2.702667E-6   -2.756204E-5   2.769424E-5   -1.743996E+2   -8.439962E+1   
4.338571E+3   1.299853E+2   1.299853E+2   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   -1.991830E-2   2.668040E-2   -2.969108E-5   -2.710698E-6   2.710698E-6   -2.969108E-5   2.981456E-5   -1.747835E+2   -8.478354E+1   
4.360588E+3   1.299694E+2   1.299694E+2   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   -2.176674E-2   2.783425E-2   -3.158537E-5   -2.097885E-6   2.097885E-6   -3.158537E-5   3.165496E-5   -1.762000E+2   -8.620002E+1   
4.382615E+3   1.300206E+2   1.300206E+2   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   -2.219134E-2   2.868252E-2   -3.240034E-5   -2.338415E-6   2.338415E-6   -3.240034E-5   3.248462E-5   -1.758720E+2   -8.587198E+1   
4.404695E+3   1.299790E+2   1.299790E+2   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.300000E+3   -1.300000E+3   -2.335594E-2   3.296566E-2   -3.590992E-5   -4.277239E-6   4.277239E-6   -3.590992E-5   3.616376E-5   -1.732075E+2   -8.320749E+1   
4.426738E+3   1.300893E+2   1.300893E+2   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   -2.416403E-2   3.267911E-2   -3.622289E-5   -3.492212E-6   3.492212E-6   -3.622289E-5   3.639084E-5   -1.744932E+2   -8.449319E+1   
4.448556E+3   1.300285E+2   1.300285E+2   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   -2.627665E-2   3.589430E-2   -3.962303E-5   -4.031651E-6   4.031651E-6   -3.962303E-5   3.982762E-5   -1.741901E+2   -8.419014E+1   
4.470647E+3   1.300135E+2   1.300135E+2   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.150000E+3   -1.150000E+3   -2.760261E-2   3.676221E-2   -4.100806E-5   -3.618348E-6   3.618348E-6   -4.100806E-5   4.116739E-5   -1.749576E+2   -8.495756E+1   
4.492662E+3   1.300568E+2   1.300568E+2   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.100000E+3   -1.100000E+3   -2.893869E-2   3.858977E-2   -4.302436E-5   -3.824949E-6   3.824949E-6   -4.302436E-5   4.319405E-5   -1.749197E+2   -8.491965E+1   
4.514743E+3   1.300073E+2   1.300073E+2   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.050000E+3   -1.050000E+3   -2.819441E-2   4.013235E-2   -4.356887E-5   -5.383932E-6   5.383932E-6   -4.356887E-5   4.390027E-5   -1.729555E+2   -8.295551E+1   
4.536761E+3   1.300420E+2   1.300420E+2   -1.000000E+3   -1.000000E+3   9.000000E+1   -1.000000E+3   -1.000000E+3   -2.926389E-2   4.171814E-2   -4.526289E-5   -5.629663E-6   5.629663E-6   -4.526289E-5   4.561165E-5   -1.729101E+2   -8.291013E+1   
4.558689E+3   1.300547E+2   1.300547E+2   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   -3.124883E-2   4.301742E-2   -4.733628E-5   -5.010967E-6   5.010967E-6   -4.733628E-5   4.760077E-5   -1.739572E+2   -8.395724E+1   
4.580413E+3   1.300497E+2   1.300497E+2   -9.000000E+2   -9.000000E+2   9.000000E+1   -8.990000E+2   -8.990000E+2   -3.271562E-2   4.446366E-2   -4.918503E-5   -4.871598E-6   4.871598E-6   -4.918503E-5   4.942570E-5   -1.743435E+2   -8.434351E+1   
4.602356E+3   1.300034E+2   1.300034E+2   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   -3.312366E-2   4.652377E-2   -5.077904E-5   -5.916638E-6   5.916638E-6   -5.077904E-5   5.112257E-5   -1.733540E+2   -8.335402E+1   
4.623989E+3   1.300498E+2   1.300498E+2   -8.000000E+2   -8.000000E+2   9.000000E+1   -8.000000E+2   -8.000000E+2   -3.392345E-2   4.711256E-2   -5.165697E-5   -5.710023E-6   5.710023E-6   -5.165697E-5   5.197160E-5   -1.736923E+2   -8.369229E+1   
4.645632E+3   1.300219E+2   1.300219E+2   -7.500000E+2   -7.500000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   -3.453429E-2   5.003912E-2   -5.394066E-5   -7.171532E-6   7.171532E-6   -5.394066E-5   5.441531E-5   -1.724268E+2   -8.242681E+1   
4.667580E+3   1.300093E+2   1.300093E+2   -7.010000E+2   -7.010000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   -3.599769E-2   5.088406E-2   -5.539571E-5   -6.641550E-6   6.641550E-6   -5.539571E-5   5.579243E-5   -1.731633E+2   -8.316328E+1   
4.689567E+3   1.300101E+2   1.300101E+2   -6.510000E+2   -6.510000E+2   9.000000E+1   -6.500000E+2   -6.500000E+2   -3.684015E-2   5.267235E-2   -5.708124E-5   -7.187576E-6   7.187576E-6   -5.708124E-5   5.753199E-5   -1.728232E+2   -8.282318E+1   
4.711295E+3   1.300347E+2   1.300347E+2   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   -3.834710E-2   5.379184E-2   -5.874203E-5   -6.804883E-6   6.804883E-6   -5.874203E-5   5.913487E-5   -1.733921E+2   -8.339211E+1   
4.733228E+3   1.300090E+2   1.300090E+2   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   -3.972029E-2   5.520615E-2   -6.051212E-5   -6.713856E-6   6.713856E-6   -6.051212E-5   6.088343E-5   -1.736689E+2   -8.366889E+1   
4.754872E+3   1.300852E+2   1.300852E+2   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   -4.142671E-2   5.738071E-2   -6.298337E-5   -6.873406E-6   6.873406E-6   -6.298337E-5   6.335731E-5   -1.737719E+2   -8.377193E+1   
4.776582E+3   1.300186E+2   1.300186E+2   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   -4.231425E-2   5.805594E-2   -6.397186E-5   -6.658403E-6   6.658403E-6   -6.397186E-5   6.431745E-5   -1.740579E+2   -8.405786E+1   
4.798252E+3   1.300449E+2   1.300449E+2   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   -4.221423E-2   6.041240E-2   -6.544477E-5   -8.272968E-6   8.272968E-6   -6.544477E-5   6.596560E-5   -1.727954E+2   -8.279537E+1   
4.819963E+3   1.300029E+2   1.300029E+2   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   -4.375157E-2   6.142237E-2   -6.705300E-5   -7.796193E-6   7.796193E-6   -6.705300E-5   6.750471E-5   -1.733680E+2   -8.336805E+1   
4.841677E+3   1.299943E+2   1.299943E+2   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   -4.515518E-2   6.330363E-2   -6.914603E-5   -7.987954E-6   7.987954E-6   -6.914603E-5   6.960590E-5   -1.734102E+2   -8.341023E+1   
4.863374E+3   1.300414E+2   1.300414E+2   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   -4.528004E-2   6.540914E-2   -7.059452E-5   -9.272129E-6   9.272129E-6   -7.059452E-5   7.120083E-5   -1.725174E+2   -8.251741E+1   
4.884995E+3   1.300535E+2   1.300535E+2   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   -4.588781E-2   6.707963E-2   -7.205824E-5   -9.914719E-6   9.914719E-6   -7.205824E-5   7.273714E-5   -1.721657E+2   -8.216569E+1   
4.906631E+3   1.299925E+2   1.299925E+2   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   -4.781882E-2   6.818745E-2   -7.397360E-5   -9.210743E-6   9.210743E-6   -7.397360E-5   7.454483E-5   -1.729024E+2   -8.290241E+1   
4.928312E+3   1.300582E+2   1.300582E+2   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   -4.875763E-2   6.951066E-2   -7.541580E-5   -9.381444E-6   9.381444E-6   -7.541580E-5   7.599707E-5   -1.729090E+2   -8.290905E+1   
4.949835E+3   1.300981E+2   1.300981E+2   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   -4.956971E-2   7.133821E-2   -7.710814E-5   -9.975612E-6   9.975612E-6   -7.710814E-5   7.775074E-5   -1.726285E+2   -8.262849E+1   
4.982870E+3   1.300041E+2   1.300041E+2   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   -4.990351E-2   7.075285E-2   -7.693327E-5   -9.346030E-6   9.346030E-6   -7.693327E-5   7.749888E-5   -1.730735E+2   -8.307352E+1   
5.005064E+3   1.300117E+2   1.300117E+2   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   -4.990290E-2   7.027363E-2   -7.662078E-5   -9.033181E-6   9.033181E-6   -7.662078E-5   7.715142E-5   -1.732762E+2   -8.327617E+1   
5.027332E+3   1.299785E+2   1.299785E+2   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   -5.032536E-2   7.049853E-2   -7.702844E-5   -8.867743E-6   8.867743E-6   -7.702844E-5   7.753720E-5   -1.734328E+2   -8.343285E+1   
5.049613E+3   1.300253E+2   1.300253E+2   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   -5.073430E-2   7.087035E-2   -7.752343E-5   -8.808367E-6   8.808367E-6   -7.752343E-5   7.802223E-5   -1.735177E+2   -8.351774E+1   
5.071864E+3   1.300300E+2   1.300300E+2   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   -4.907454E-2   7.174994E-2   -7.707015E-5   -1.061103E-5   1.061103E-5   -7.707015E-5   7.779718E-5   -1.721608E+2   -8.216079E+1   
5.094129E+3   1.300299E+2   1.300299E+2   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   -4.925555E-2   7.199536E-2   -7.734190E-5   -1.063760E-5   1.063760E-5   -7.734190E-5   7.807002E-5   -1.721687E+2   -8.216868E+1   
5.116364E+3   1.300093E+2   1.300093E+2   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   -5.098315E-2   7.121794E-2   -7.790366E-5   -8.851560E-6   8.851560E-6   -7.790366E-5   7.840491E-5   -1.735177E+2   -8.351775E+1   
5.138636E+3   1.300539E+2   1.300539E+2   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   -4.973081E-2   7.109951E-2   -7.705227E-5   -9.700401E-6   9.700401E-6   -7.705227E-5   7.766048E-5   -1.728246E+2   -8.282457E+1   
5.160918E+3   1.300252E+2   1.300252E+2   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   -5.012348E-2   7.150143E-2   -7.755680E-5   -9.672727E-6   9.672727E-6   -7.755680E-5   7.815766E-5   -1.728909E+2   -8.289089E+1   
5.183238E+3   1.299773E+2   1.299773E+2   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   -4.919666E-2   7.072645E-2   -7.647906E-5   -9.851582E-6   9.851582E-6   -7.647906E-5   7.711096E-5   -1.726599E+2   -8.265992E+1   
5.205431E+3   1.300443E+2   1.300443E+2   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   -5.098068E-2   7.189228E-2   -7.834132E-5   -9.294244E-6   9.294244E-6   -7.834132E-5   7.889072E-5   -1.732342E+2   -8.323418E+1   
5.227705E+3   1.299634E+2   1.299634E+2   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   -4.984246E-2   7.247366E-2   -7.801627E-5   -1.051620E-5   1.051620E-5   -7.801627E-5   7.872185E-5   -1.723231E+2   -8.232309E+1   
5.249969E+3   1.300297E+2   1.300297E+2   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   -4.941695E-2   7.235798E-2   -7.767786E-5   -1.075530E-5   1.075530E-5   -7.767786E-5   7.841891E-5   -1.721169E+2   -8.211693E+1   
5.272216E+3   1.299928E+2   1.299928E+2   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   -4.966175E-2   7.225673E-2   -7.776326E-5   -1.050804E-5   1.050804E-5   -7.776326E-5   7.847002E-5   -1.723043E+2   -8.230432E+1   
5.294489E+3   1.300485E+2   1.300485E+2   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   -5.090859E-2   7.180485E-2   -7.823981E-5   -9.290406E-6   9.290406E-6   -7.823981E-5   7.878946E-5   -1.732283E+2   -8.322825E+1   
5.316732E+3   1.300433E+2   1.300433E+2   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   -4.987928E-2   7.252489E-2   -7.807239E-5   -1.052246E-5   1.052246E-5   -7.807239E-5   7.877830E-5   -1.723240E+2   -8.232403E+1   
5.338923E+3   1.300138E+2   1.300138E+2   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   -4.969857E-2   7.293445E-2   -7.822742E-5   -1.092388E-5   1.092388E-5   -7.822742E-5   7.898645E-5   -1.720505E+2   -8.205047E+1   
5.361165E+3   1.299848E+2   1.299848E+2   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   -5.023304E-2   7.209783E-2   -7.801297E-5   -9.981610E-6   9.981610E-6   -7.801297E-5   7.864894E-5   -1.727087E+2   -8.270873E+1   
5.383417E+3   1.299687E+2   1.299687E+2   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   -5.048459E-2   7.272461E-2   -7.857671E-5   -1.020533E-5   1.020533E-5   -7.857671E-5   7.923665E-5   -1.726000E+2   -8.260001E+1   
5.405496E+3   1.300443E+2   1.300443E+2   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   -4.914727E-2   7.246690E-2   -7.758207E-5   -1.102597E-5   1.102597E-5   -7.758207E-5   7.836166E-5   -1.719113E+2   -8.191129E+1   
5.427543E+3   1.300123E+2   1.300123E+2   -8.000000E+0   -8.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   -5.061987E-2   7.267123E-2   -7.862557E-5   -1.007037E-5   1.007037E-5   -7.862557E-5   7.926786E-5   -1.727013E+2   -8.270129E+1   
5.449620E+3   1.299622E+2   1.299622E+2   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   -5.003205E-2   7.281511E-2   -7.835586E-5   -1.059920E-5   1.059920E-5   -7.835586E-5   7.906949E-5   -1.722964E+2   -8.229636E+1   
5.471646E+3   1.300457E+2   1.300457E+2   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   -5.017196E-2   7.282985E-2   -7.845196E-5   -1.050536E-5   1.050536E-5   -7.845196E-5   7.915221E-5   -1.723730E+2   -8.237300E+1   
5.493732E+3   1.300861E+2   1.300861E+2   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   -4.999433E-2   7.200764E-2   -7.780665E-5   -1.009920E-5   1.009920E-5   -7.780665E-5   7.845934E-5   -1.726044E+2   -8.260443E+1   
5.515709E+3   1.300189E+2   1.300189E+2   0.000000E+0   0.000000E+0   9.000000E+1   0.000000E+0   0.000000E+0   -5.028946E-2   7.376034E-2   -7.913062E-5   -1.102678E-5   1.102678E-5   -7.913062E-5   7.989522E-5   -1.720670E+2   -8.206697E+1   
5.537693E+3   1.300083E+2   1.300083E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   -5.102363E-2   7.369437E-2   -7.954156E-5   -1.044064E-5   1.044064E-5   -7.954156E-5   8.022385E-5   -1.725221E+2   -8.252210E+1   
5.559222E+3   1.299586E+2   1.299586E+2   3.000000E+0   3.000000E+0   9.000000E+1   3.000000E+0   3.000000E+0   -4.977622E-2   7.331118E-2   -7.852078E-5   -1.111275E-5   1.111275E-5   -7.852078E-5   7.930326E-5   -1.719446E+2   -8.194465E+1   
5.580880E+3   1.300412E+2   1.300412E+2   5.000000E+0   5.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   -4.955347E-2   7.382601E-2   -7.871837E-5   -1.161408E-5   1.161408E-5   -7.871837E-5   7.957052E-5   -1.716072E+2   -8.160715E+1   
5.602595E+3   1.300436E+2   1.300436E+2   6.000000E+0   6.000000E+0   9.000000E+1   8.000000E+0   8.000000E+0   -5.226554E-2   7.295194E-2   -7.982583E-5   -9.036705E-6   9.036705E-6   -7.982583E-5   8.033570E-5   -1.735413E+2   -8.354131E+1   
5.624184E+3   1.299533E+2   1.299533E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   -5.081779E-2   7.340232E-2   -7.922408E-5   -1.040195E-5   1.040195E-5   -7.922408E-5   7.990404E-5   -1.725200E+2   -8.251998E+1   
5.646043E+3   1.299119E+2   1.299119E+2   1.000000E+1   1.000000E+1   9.000000E+1   1.100000E+1   1.100000E+1   -5.075087E-2   7.285039E-2   -7.882325E-5   -1.009060E-5   1.009060E-5   -7.882325E-5   7.946650E-5   -1.727049E+2   -8.270493E+1   
5.667952E+3   1.300109E+2   1.300109E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   -5.027137E-2   7.297648E-2   -7.860892E-5   -1.052769E-5   1.052769E-5   -7.860892E-5   7.931074E-5   -1.723721E+2   -8.237206E+1   
5.689849E+3   1.299810E+2   1.299810E+2   1.500000E+1   1.500000E+1   9.000000E+1   1.600000E+1   1.600000E+1   -5.109328E-2   7.323419E-2   -7.928491E-5   -1.008827E-5   1.008827E-5   -7.928491E-5   7.992415E-5   -1.727486E+2   -8.274861E+1   
5.711884E+3   1.299510E+2   1.299510E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   -5.151297E-2   7.275313E-2   -7.923107E-5   -9.463347E-6   9.463347E-6   -7.923107E-5   7.979422E-5   -1.731889E+2   -8.318887E+1   
5.733727E+3   1.299372E+2   1.299372E+2   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   -4.942706E-2   7.419354E-2   -7.887959E-5   -1.194785E-5   1.194785E-5   -7.887959E-5   7.977932E-5   -1.713869E+2   -8.138691E+1   
5.755660E+3   1.300161E+2   1.300161E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   -5.099202E-2   7.404628E-2   -7.975121E-5   -1.069408E-5   1.069408E-5   -7.975121E-5   8.046501E-5   -1.723626E+2   -8.236259E+1   
5.777522E+3   1.300755E+2   1.300755E+2   2.200000E+1   2.200000E+1   9.000000E+1   2.300000E+1   2.300000E+1   -4.995873E-2   7.381679E-2   -7.896291E-5   -1.130830E-5   1.130830E-5   -7.896291E-5   7.976854E-5   -1.718501E+2   -8.185007E+1   
5.799395E+3   1.300368E+2   1.300368E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   -5.082054E-2   7.257736E-2   -7.868850E-5   -9.860578E-6   9.860578E-6   -7.868850E-5   7.930392E-5   -1.728574E+2   -8.285741E+1   
5.821276E+3   1.300008E+2   1.300008E+2   2.600000E+1   2.600000E+1   9.000000E+1   2.700000E+1   2.700000E+1   -5.084356E-2   7.297648E-2   -7.896268E-5   -1.010448E-5   1.010448E-5   -7.896268E-5   7.960656E-5   -1.727078E+2   -8.270776E+1   
5.843151E+3   1.299730E+2   1.299730E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   -5.036340E-2   7.289426E-2   -7.861227E-5   -1.040587E-5   1.040587E-5   -7.861227E-5   7.929799E-5   -1.724596E+2   -8.245962E+1   
5.865034E+3   1.300271E+2   1.300271E+2   3.100000E+1   3.100000E+1   9.000000E+1   3.100000E+1   3.100000E+1   -5.062049E-2   7.482123E-2   -8.002623E-5   -1.147552E-5   1.147552E-5   -8.002623E-5   8.084482E-5   -1.718396E+2   -8.183959E+1   
5.887163E+3   1.300266E+2   1.300266E+2   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   -5.117549E-2   7.382813E-2   -7.972256E-5   -1.041576E-5   1.041576E-5   -7.972256E-5   8.040009E-5   -1.725565E+2   -8.255646E+1   
5.909103E+3   1.300849E+2   1.300849E+2   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   -5.154487E-2   7.397355E-2   -8.004564E-5   -1.023763E-5   1.023763E-5   -8.004564E-5   8.069767E-5   -1.727116E+2   -8.271158E+1   
5.931030E+3   1.300385E+2   1.300385E+2   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   -5.094908E-2   7.311115E-2   -7.911562E-5   -1.011448E-5   1.011448E-5   -7.911562E-5   7.975954E-5   -1.727146E+2   -8.271458E+1   
5.952998E+3   1.300073E+2   1.300073E+2   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   -5.139363E-2   7.319124E-2   -7.944263E-5   -9.838046E-6   9.838046E-6   -7.944263E-5   8.004947E-5   -1.729405E+2   -8.294053E+1   
5.974873E+3   1.300865E+2   1.300865E+2   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   -5.074202E-2   7.435090E-2   -7.979504E-5   -1.107815E-5   1.107815E-5   -7.979504E-5   8.056037E-5   -1.720960E+2   -8.209600E+1   
5.996797E+3   1.300372E+2   1.300372E+2   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   -5.147554E-2   7.444572E-2   -8.031030E-5   -1.059760E-5   1.059760E-5   -8.031030E-5   8.100650E-5   -1.724828E+2   -8.248279E+1   
6.018654E+3   1.300224E+2   1.300224E+2   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   -5.195076E-2   7.401039E-2   -8.032057E-5   -9.961504E-6   9.961504E-6   -8.032057E-5   8.093594E-5   -1.729302E+2   -8.293017E+1   
6.040536E+3   1.300126E+2   1.300126E+2   4.600000E+1   4.600000E+1   9.000000E+1   4.800000E+1   4.800000E+1   -5.095092E-2   7.347563E-2   -7.935414E-5   -1.035141E-5   1.035141E-5   -7.935414E-5   8.002644E-5   -1.725680E+2   -8.256797E+1   
6.062418E+3   1.300626E+2   1.300626E+2   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   -4.943011E-2   7.513752E-2   -7.949628E-5   -1.256274E-5   1.256274E-5   -7.949628E-5   8.048280E-5   -1.710198E+2   -8.101985E+1   
6.096316E+3   1.300312E+2   1.300312E+2   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   -5.290798E-2   7.622174E-2   -8.235260E-5   -1.069923E-5   1.069923E-5   -8.235260E-5   8.304471E-5   -1.725976E+2   -8.259761E+1   
6.119106E+3   1.299461E+2   1.299461E+2   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   -5.258982E-2   7.726974E-2   -8.283845E-5   -1.161971E-5   1.161971E-5   -8.283845E-5   8.364942E-5   -1.720152E+2   -8.201525E+1   
6.141320E+3   1.300748E+2   1.300748E+2   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   -5.407746E-2   7.893286E-2   -8.484135E-5   -1.160671E-5   1.160671E-5   -8.484135E-5   8.563160E-5   -1.722100E+2   -8.221002E+1   
6.163476E+3   1.299948E+2   1.299948E+2   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   -5.551876E-2   8.106323E-2   -8.711992E-5   -1.193345E-5   1.193345E-5   -8.711992E-5   8.793343E-5   -1.722003E+2   -8.220032E+1   
6.186075E+3   1.300312E+2   1.300312E+2   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   -5.647443E-2   8.109975E-2   -8.773454E-5   -1.125048E-5   1.125048E-5   -8.773454E-5   8.845294E-5   -1.726927E+2   -8.269266E+1   
6.208475E+3   1.300201E+2   1.300201E+2   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   -5.767889E-2   8.435265E-2   -9.059778E-5   -1.248628E-5   1.248628E-5   -9.059778E-5   9.145416E-5   -1.721529E+2   -8.215287E+1   
6.230801E+3   1.300063E+2   1.300063E+2   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   -5.872321E-2   8.497393E-2   -9.164806E-5   -1.212004E-5   1.212004E-5   -9.164806E-5   9.244599E-5   -1.724666E+2   -8.246661E+1   
6.253680E+3   1.300248E+2   1.300248E+2   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   -6.013691E-2   8.695334E-2   -9.381124E-5   -1.236851E-5   1.236851E-5   -9.381124E-5   9.462308E-5   -1.724892E+2   -8.248918E+1   
6.275801E+3   1.299431E+2   1.299431E+2   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   -6.157976E-2   8.856278E-2   -9.575149E-5   -1.235355E-5   1.235355E-5   -9.575149E-5   9.654511E-5   -1.726485E+2   -8.264849E+1   
6.298410E+3   1.300525E+2   1.300525E+2   5.480000E+2   5.480000E+2   9.000000E+1   5.480000E+2   5.480000E+2   -6.258512E-2   8.996148E-2   -9.728401E-5   -1.252437E-5   1.252437E-5   -9.728401E-5   9.808689E-5   -1.726641E+2   -8.266407E+1   
6.321770E+3   1.301263E+2   1.301263E+2   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   -6.231791E-2   9.079842E-2   -9.766390E-5   -1.326918E-5   1.326918E-5   -9.766390E-5   9.856119E-5   -1.722628E+2   -8.226284E+1   
6.344460E+3   1.300345E+2   1.300345E+2   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   -6.453324E-2   9.278038E-2   -1.003243E-4   -1.292640E-5   1.292640E-5   -1.003243E-4   1.011537E-4   -1.726581E+2   -8.265811E+1   
6.367334E+3   1.299553E+2   1.299553E+2   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   -6.554719E-2   9.427545E-2   -1.019249E-4   -1.315389E-5   1.315389E-5   -1.019249E-4   1.027702E-4   -1.726464E+2   -8.264636E+1   
6.390715E+3   1.300514E+2   1.300514E+2   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   -6.577638E-2   9.641757E-2   -1.034618E-4   -1.438483E-5   1.438483E-5   -1.034618E-4   1.044570E-4   -1.720846E+2   -8.208462E+1   
6.413394E+3   1.300204E+2   1.300204E+2   7.970000E+2   7.970000E+2   9.000000E+1   7.980000E+2   7.980000E+2   -6.758554E-2   9.794821E-2   -1.055772E-4   -1.404740E-5   1.404740E-5   -1.055772E-4   1.065076E-4   -1.724211E+2   -8.242111E+1   
6.436034E+3   1.299738E+2   1.299738E+2   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   -6.847063E-2   9.938861E-2   -1.070625E-4   -1.433446E-5   1.433446E-5   -1.070625E-4   1.080178E-4   -1.723741E+2   -8.237409E+1   
6.459375E+3   1.299313E+2   1.299313E+2   8.980000E+2   8.980000E+2   9.000000E+1   8.980000E+2   8.980000E+2   -6.804173E-2   1.006756E-1   -1.076355E-4   -1.549308E-5   1.549308E-5   -1.076355E-4   1.087448E-4   -1.718091E+2   -8.180909E+1   
6.481925E+3   1.300838E+2   1.300838E+2   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   -7.072587E-2   1.013880E-1   -1.097590E-4   -1.397355E-5   1.397355E-5   -1.097590E-4   1.106449E-4   -1.727446E+2   -8.274463E+1   
6.504556E+3   1.300254E+2   1.300254E+2   9.980000E+2   9.980000E+2   9.000000E+1   9.980000E+2   9.980000E+2   -7.110996E-2   1.034496E-1   -1.113392E-4   -1.503731E-5   1.503731E-5   -1.113392E-4   1.123500E-4   -1.723083E+2   -8.230825E+1   
6.528030E+3   1.300657E+2   1.300657E+2   1.048000E+3   1.048000E+3   9.000000E+1   1.048000E+3   1.048000E+3   -7.178799E-2   1.047062E-1   -1.125768E-4   -1.535736E-5   1.535736E-5   -1.125768E-4   1.136194E-4   -1.722318E+2   -8.223184E+1   
6.550782E+3   1.299497E+2   1.299497E+2   1.098000E+3   1.098000E+3   9.000000E+1   1.098000E+3   1.098000E+3   -7.354744E-2   1.071321E-1   -1.152444E-4   -1.564194E-5   1.564194E-5   -1.152444E-4   1.163011E-4   -1.722706E+2   -8.227057E+1   
6.573535E+3   1.300369E+2   1.300369E+2   1.148000E+3   1.148000E+3   9.000000E+1   1.149000E+3   1.149000E+3   -7.434879E-2   1.082374E-1   -1.164598E-4   -1.577190E-5   1.577190E-5   -1.164598E-4   1.175229E-4   -1.722875E+2   -8.228748E+1   
6.596792E+3   1.299945E+2   1.299945E+2   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   -7.486206E-2   1.097702E-1   -1.177754E-4   -1.639434E-5   1.639434E-5   -1.177754E-4   1.189109E-4   -1.720753E+2   -8.207535E+1   
6.619619E+3   1.300510E+2   1.300510E+2   1.248000E+3   1.248000E+3   9.000000E+1   1.248000E+3   1.248000E+3   -7.556459E-2   1.103387E-1   -1.185800E-4   -1.624639E-5   1.624639E-5   -1.185800E-4   1.196877E-4   -1.721986E+2   -8.219860E+1   
6.642670E+3   1.300738E+2   1.300738E+2   1.297000E+3   1.297000E+3   9.000000E+1   1.299000E+3   1.299000E+3   -7.715930E-2   1.124285E-1   -1.209270E-4   -1.643318E-5   1.643318E-5   -1.209270E-4   1.220385E-4   -1.722613E+2   -8.226129E+1   
6.666272E+3   1.299963E+2   1.299963E+2   1.348000E+3   1.348000E+3   9.000000E+1   1.348000E+3   1.348000E+3   -7.808643E-2   1.137263E-1   -1.223454E-4   -1.659587E-5   1.659587E-5   -1.223454E-4   1.234658E-4   -1.722751E+2   -8.227511E+1   
6.688806E+3   1.300986E+2   1.300986E+2   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   -7.852728E-2   1.150909E-1   -1.235067E-4   -1.716195E-5   1.716195E-5   -1.235067E-4   1.246934E-4   -1.720891E+2   -8.208909E+1   
6.711431E+3   1.300707E+2   1.300707E+2   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   -7.975018E-2   1.162395E-1   -1.250109E-4   -1.700841E-5   1.700841E-5   -1.250109E-4   1.261626E-4   -1.722522E+2   -8.225217E+1   
6.734206E+3   1.300213E+2   1.300213E+2   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   -7.985047E-2   1.179582E-1   -1.261922E-4   -1.805782E-5   1.805782E-5   -1.261922E-4   1.274777E-4   -1.718564E+2   -8.185639E+1   
6.756783E+3   1.300584E+2   1.300584E+2   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   -8.143169E-2   1.190252E-1   -1.278647E-4   -1.758590E-5   1.758590E-5   -1.278647E-4   1.290684E-4   -1.721689E+2   -8.216894E+1   
6.779380E+3   1.300457E+2   1.300457E+2   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   -8.304020E-2   1.209040E-1   -1.300828E-4   -1.762450E-5   1.762450E-5   -1.300828E-4   1.312713E-4   -1.722842E+2   -8.228416E+1   
6.802385E+3   1.300000E+2   1.300000E+2   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   -8.285552E-2   1.221471E-1   -1.307783E-4   -1.857381E-5   1.857381E-5   -1.307783E-4   1.320907E-4   -1.719166E+2   -8.191662E+1   
6.824963E+3   1.300489E+2   1.300489E+2   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   -8.476591E-2   1.243459E-1   -1.333914E-4   -1.859833E-5   1.859833E-5   -1.333914E-4   1.346817E-4   -1.720626E+2   -8.206261E+1   
6.847484E+3   1.300366E+2   1.300366E+2   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   -8.487912E-2   1.251092E-1   -1.339585E-4   -1.901363E-5   1.901363E-5   -1.339585E-4   1.353012E-4   -1.719216E+2   -8.192159E+1   
6.870258E+3   1.301160E+2   1.301160E+2   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   -8.676223E-2   1.277056E-1   -1.368138E-4   -1.931826E-5   1.931826E-5   -1.368138E-4   1.381709E-4   -1.719629E+2   -8.196290E+1   
6.892821E+3   1.300675E+2   1.300675E+2   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   -8.812068E-2   1.293144E-1   -1.387014E-4   -1.936530E-5   1.936530E-5   -1.387014E-4   1.400468E-4   -1.720518E+2   -8.205182E+1   
6.915352E+3   1.299745E+2   1.299745E+2   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   -8.997036E-2   1.311162E-1   -1.410185E-4   -1.917518E-5   1.917518E-5   -1.410185E-4   1.423162E-4   -1.722566E+2   -8.225662E+1   
6.938136E+3   1.299538E+2   1.299538E+2   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   -9.136513E-2   1.337101E-1   -1.435702E-4   -1.983941E-5   1.983941E-5   -1.435702E-4   1.449345E-4   -1.721323E+2   -8.213234E+1   
6.960703E+3   1.299635E+2   1.299635E+2   1.999000E+3   1.999000E+3   9.000000E+1   1.999000E+3   1.999000E+3   -9.043025E-2   1.349928E-1   -1.438276E-4   -2.136948E-5   2.136948E-5   -1.438276E-4   1.454064E-4   -1.715490E+2   -8.154899E+1   
6.998601E+3   1.300123E+2   1.300123E+2   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   -1.045750E-1   1.516664E-1   -1.634318E-4   -2.180829E-5   2.180829E-5   -1.634318E-4   1.648805E-4   -1.723994E+2   -8.239937E+1   
7.025538E+3   1.300105E+2   1.300105E+2   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   -1.162954E-1   1.691759E-1   -1.820817E-4   -2.458680E-5   2.458680E-5   -1.820817E-4   1.837342E-4   -1.723098E+2   -8.230977E+1   
7.051468E+3   1.300732E+2   1.300732E+2   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -1.252721E-1   1.850025E-1   -1.979393E-4   -2.829429E-5   2.829429E-5   -1.979393E-4   1.999513E-4   -1.718650E+2   -8.186500E+1   
7.077158E+3   1.299688E+2   1.299688E+2   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -1.319994E-1   1.976703E-1   -2.103488E-4   -3.160041E-5   3.160041E-5   -2.103488E-4   2.127092E-4   -1.714564E+2   -8.145643E+1   
7.103756E+3   1.299263E+2   1.299263E+2   4.498000E+3   4.498000E+3   9.000000E+1   4.499000E+3   4.499000E+3   -1.362129E-1   2.032920E-1   -2.166151E-4   -3.215926E-5   3.215926E-5   -2.166151E-4   2.189894E-4   -1.715554E+2   -8.155540E+1   
7.129721E+3   1.299750E+2   1.299750E+2   4.998000E+3   4.998000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -1.250945E-1   1.951598E-1   -2.044448E-4   -3.506624E-5   3.506624E-5   -2.044448E-4   2.074303E-4   -1.702674E+2   -8.026737E+1   
7.155369E+3   1.300407E+2   1.300407E+2   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -1.122129E-1   1.783997E-1   -1.855650E-4   -3.363654E-5   3.363654E-5   -1.855650E-4   1.885890E-4   -1.697258E+2   -7.972581E+1   
7.181818E+3   1.299989E+2   1.299989E+2   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -9.662557E-2   1.624327E-1   -1.655291E-4   -3.472661E-5   3.472661E-5   -1.655291E-4   1.691326E-4   -1.681517E+2   -7.815166E+1   
7.207746E+3   1.300702E+2   1.300702E+2   6.498000E+3   6.498000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -8.415693E-2   1.494931E-1   -1.493930E-4   -3.548926E-5   3.548926E-5   -1.493930E-4   1.535505E-4   -1.666367E+2   -7.663672E+1   
7.233947E+3   1.299914E+2   1.299914E+2   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -7.989559E-2   1.513381E-1   -1.479601E-4   -3.984732E-5   3.984732E-5   -1.479601E-4   1.532318E-4   -1.649272E+2   -7.492721E+1   
7.259638E+3   1.299976E+2   1.299976E+2   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -8.480119E-2   1.557970E-1   -1.538970E-4   -3.913412E-5   3.913412E-5   -1.538970E-4   1.587947E-4   -1.657328E+2   -7.573278E+1   
7.285062E+3   1.300538E+2   1.300538E+2   7.999000E+3   7.999000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -9.639543E-2   1.719435E-1   -1.715812E-4   -4.111476E-5   4.111476E-5   -1.715812E-4   1.764384E-4   -1.665247E+2   -7.652470E+1   
7.311491E+3   1.300339E+2   1.300339E+2   8.498000E+3   8.498000E+3   9.000000E+1   8.499000E+3   8.499000E+3   -1.017800E-1   1.829081E-1   -1.820513E-4   -4.430046E-5   4.430046E-5   -1.820513E-4   1.873638E-4   -1.663234E+2   -7.632343E+1   
7.337887E+3   1.299991E+2   1.299991E+2   8.998000E+3   8.998000E+3   9.000000E+1   8.999000E+3   8.999000E+3   -1.115342E-1   1.998409E-1   -1.991099E-4   -4.815615E-5   4.815615E-5   -1.991099E-4   2.048506E-4   -1.664037E+2   -7.640370E+1   
7.364289E+3   1.300149E+2   1.300149E+2   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -1.189902E-1   2.137361E-1   -2.127694E-4   -5.172579E-5   5.172579E-5   -2.127694E-4   2.189666E-4   -1.663360E+2   -7.633605E+1   
7.389684E+3   1.299925E+2   1.299925E+2   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -1.341755E-1   2.338065E-1   -2.352293E-4   -5.361572E-5   5.361572E-5   -2.352293E-4   2.412622E-4   -1.671600E+2   -7.715995E+1   
@@END Data.
@Time at end of measurement: 17:36:08
@NO Instrument  Changes.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -9499.000      -9999.000      250.000        Coercive Field: Field at which M//H changes sign
Ms  emu                                 3.139E-4       -3.002E-4      3.070E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -7.913E-5      1.435E-4       1.113E-4       Remanent Magnetization: M at H=0        
S                                       0.252          0.478          0.365          Squareness: Mr/Ms                       
S*                                      1.318          1.195          1.256          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
