@Filename: c:\vsm-lv\Will\data\AJA335e-FePtFeRh_1030nm_Tann_6\AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_110deg.VHD
@Measurement Controlfilename: C:\vsm-lv\Will\Recipes\10kOe OoP loop 110deg.VHC
@Signal Manipulation filename: c:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA335e-FePtFeRh_1030nm_Tann_6
@Date: 08 November 2019    (2019-08-11)
@Time: 10:52:16
@Test ID: AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_110deg
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 90.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Sample Temperature to 110.0942 [degC] and wait 60.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Applied Field to 9999.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 3:      Set Auto Range Signal to 12.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 5
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 5.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 10000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To: 50.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: 50.0000 [Oe] To: -50.0000 [Oe] Min Stepsize/Sweeprate =  2.0000 [Oe] Max Stepsize/Sweeprate =  2.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -50.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -10000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 4 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 20 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.706
@Y Coils Correction Factor: 0.964
@Sample Shape Correction Factor: 0.919
@Coil Angle Alpha: 42.300
@Coil Angle Beta: -47.320
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
15000.000000   1.000000
15249.000000   1.000524
15499.000000   1.000702
15750.000000   1.001233
16000.000000   1.001406
16250.000000   1.001585
16499.000000   1.001758
16749.000000   1.001937
16999.000000   1.002110
17249.000000   1.001937
17499.000000   1.002289
17749.000000   1.002289
17999.000000   1.002289
18249.000000   1.002462
18499.000000   1.002462
18748.000000   1.002462
18999.000000   1.002462
19249.000000   1.002462
19499.000000   1.002642
19749.000000   1.002642
19999.000000   1.002462
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = No
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 25 October 2019  12:02:56
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 5
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 10:52:16
@@Data
New Section: Section 0: 
3.211900E+1   1.100950E+2   1.100950E+2   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -2.131127E-1   2.984384E-1   -3.261261E-4   -3.748582E-5   3.748582E-5   -3.261261E-4   3.282734E-4   -1.734430E+2   -8.344304E+1   
5.695400E+1   1.100253E+2   1.100253E+2   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -1.939664E-1   2.762141E-1   -2.998144E-4   -3.711741E-5   3.711741E-5   -2.998144E-4   3.021032E-4   -1.729426E+2   -8.294262E+1   
8.208400E+1   1.100851E+2   1.100851E+2   8.998000E+3   8.998000E+3   9.000000E+1   8.998000E+3   8.998000E+3   -1.734333E-1   2.501733E-1   -2.701598E-4   -3.527960E-5   3.527960E-5   -2.701598E-4   2.724536E-4   -1.725600E+2   -8.255997E+1   
1.074360E+2   1.100547E+2   1.100547E+2   8.498000E+3   8.498000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -1.592479E-1   2.303625E-1   -2.484871E-4   -3.281981E-5   3.281981E-5   -2.484871E-4   2.506451E-4   -1.724760E+2   -8.247601E+1   
1.327680E+2   1.100624E+2   1.100624E+2   7.998000E+3   7.998000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -1.436744E-1   2.076601E-1   -2.240731E-4   -2.949626E-5   2.949626E-5   -2.240731E-4   2.260062E-4   -1.725009E+2   -8.250088E+1   
1.583240E+2   1.100422E+2   1.100422E+2   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -1.258455E-1   1.850931E-1   -1.983527E-4   -2.792940E-5   2.792940E-5   -1.983527E-4   2.003094E-4   -1.719851E+2   -8.198506E+1   
1.832040E+2   1.100381E+2   1.100381E+2   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -1.116444E-1   1.658147E-1   -1.770172E-4   -2.582935E-5   2.582935E-5   -1.770172E-4   1.788917E-4   -1.716983E+2   -8.169831E+1   
2.086170E+2   1.099853E+2   1.099853E+2   6.497000E+3   6.497000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -9.480655E-2   1.444242E-1   -1.526758E-4   -2.429863E-5   2.429863E-5   -1.526758E-4   1.545973E-4   -1.709571E+2   -8.095712E+1   
2.337530E+2   1.100559E+2   1.100559E+2   5.998000E+3   5.998000E+3   9.000000E+1   5.998000E+3   5.998000E+3   -8.356176E-2   1.259286E-1   -1.336778E-4   -2.052371E-5   2.052371E-5   -1.336778E-4   1.352441E-4   -1.712715E+2   -8.127147E+1   
2.593910E+2   1.100841E+2   1.100841E+2   5.498000E+3   5.498000E+3   9.000000E+1   5.498000E+3   5.498000E+3   -6.765795E-2   1.050002E-1   -1.102148E-4   -1.860422E-5   1.860422E-5   -1.102148E-4   1.117740E-4   -1.704188E+2   -8.041881E+1   
2.847880E+2   1.100144E+2   1.100144E+2   4.997000E+3   4.997000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -5.084228E-2   8.221064E-2   -8.497599E-5   -1.614247E-5   1.614247E-5   -8.497599E-5   8.649566E-5   -1.692440E+2   -7.924396E+1   
3.099260E+2   1.100146E+2   1.100146E+2   4.498000E+3   4.498000E+3   9.000000E+1   4.498000E+3   4.498000E+3   -3.707331E-2   6.365215E-2   -6.437643E-5   -1.419341E-5   1.419341E-5   -6.437643E-5   6.592251E-5   -1.675666E+2   -7.756661E+1   
3.356850E+2   1.100208E+2   1.100208E+2   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -2.000851E-2   4.126040E-2   -3.924266E-5   -1.217597E-5   1.217597E-5   -3.924266E-5   4.108821E-5   -1.627622E+2   -7.276225E+1   
3.614460E+2   1.099885E+2   1.099885E+2   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -7.872644E-3   2.167593E-2   -1.898454E-5   -8.348261E-6   8.348261E-6   -1.898454E-5   2.073900E-5   -1.562630E+2   -6.626299E+1   
3.867960E+2   1.100648E+2   1.100648E+2   2.998000E+3   2.998000E+3   9.000000E+1   2.998000E+3   2.998000E+3   9.061477E-3   1.868683E-3   4.385176E-6   -7.923842E-6   7.923842E-6   4.385176E-6   9.056326E-6   -6.103918E+1   2.896082E+1   
4.126450E+2   1.099576E+2   1.099576E+2   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   2.400604E-2   -1.962347E-2   2.762222E-5   -4.926345E-6   4.926345E-6   2.762222E-5   2.805808E-5   -1.011222E+1   7.988778E+1   
4.384880E+2   1.100373E+2   1.100373E+2   1.998000E+3   1.998000E+3   9.000000E+1   1.999000E+3   1.999000E+3   3.931749E-2   -4.002035E-2   5.037274E-5   -2.916264E-6   2.916264E-6   5.037274E-5   5.045709E-5   -3.313366E+0   8.668663E+1   
4.723690E+2   1.100256E+2   1.100256E+2   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   4.161229E-2   -4.188074E-2   5.300315E-5   -3.397293E-6   3.397293E-6   5.300315E-5   5.311191E-5   -3.667417E+0   8.633258E+1   
4.946590E+2   1.100482E+2   1.100482E+2   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   4.401267E-2   -4.432988E-2   5.608227E-5   -3.571516E-6   3.571516E-6   5.608227E-5   5.619588E-5   -3.643876E+0   8.635612E+1   
5.169780E+2   1.100815E+2   1.100815E+2   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   4.479809E-2   -4.572797E-2   5.747841E-5   -3.238400E-6   3.238400E-6   5.747841E-5   5.756957E-5   -3.224701E+0   8.677530E+1   
5.392080E+2   1.099422E+2   1.099422E+2   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   4.685731E-2   -4.894663E-2   6.084780E-5   -2.657197E-6   2.657197E-6   6.084780E-5   6.090579E-5   -2.500493E+0   8.749951E+1   
5.614420E+2   1.100069E+2   1.100069E+2   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   4.797373E-2   -5.056037E-2   6.258904E-5   -2.427922E-6   2.427922E-6   6.258904E-5   6.263611E-5   -2.221474E+0   8.777853E+1   
5.837210E+2   1.100231E+2   1.100231E+2   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   5.088554E-2   -5.251098E-2   6.565967E-5   -3.306328E-6   3.306328E-6   6.565967E-5   6.574286E-5   -2.882725E+0   8.711727E+1   
6.059460E+2   1.099879E+2   1.099879E+2   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   4.977406E-2   -5.551264E-2   6.692745E-5   -5.218395E-7   5.218395E-7   6.692745E-5   6.692948E-5   -4.467314E-1   8.955327E+1   
6.279410E+2   1.101226E+2   1.101226E+2   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   5.259105E-2   -5.634435E-2   6.921072E-5   -2.061628E-6   2.061628E-6   6.921072E-5   6.924142E-5   -1.706204E+0   8.829380E+1   
6.501790E+2   1.100378E+2   1.100378E+2   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   5.485855E-2   -5.893765E-2   7.230159E-5   -2.043313E-6   2.043313E-6   7.230159E-5   7.233045E-5   -1.618804E+0   8.838120E+1   
6.724260E+2   1.100306E+2   1.100306E+2   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   5.494536E-2   -6.077322E-2   7.355074E-5   -9.074829E-7   9.074829E-7   7.355074E-5   7.355634E-5   -7.068902E-1   8.929311E+1   
6.947070E+2   1.100370E+2   1.100370E+2   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   5.668212E-2   -6.174574E-2   7.525788E-5   -1.556242E-6   1.556242E-6   7.525788E-5   7.527397E-5   -1.184639E+0   8.881536E+1   
7.172290E+2   1.100076E+2   1.100076E+2   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   5.956874E-2   -6.510759E-2   7.923206E-5   -1.493390E-6   1.493390E-6   7.923206E-5   7.924614E-5   -1.079800E+0   8.892020E+1   
7.395350E+2   1.099982E+2   1.099982E+2   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   5.899012E-2   -6.784785E-2   8.065904E-5   7.260796E-7   -7.260796E-7   8.065904E-5   8.066231E-5   5.157534E-1   9.051575E+1   
7.617780E+2   1.099845E+2   1.099845E+2   1.297000E+3   1.297000E+3   9.000000E+1   1.299000E+3   1.299000E+3   6.095451E-2   -6.829391E-2   8.216403E-5   -4.352233E-7   4.352233E-7   8.216403E-5   8.216518E-5   -3.034932E-1   8.969651E+1   
7.840530E+2   1.100156E+2   1.100156E+2   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   6.078947E-2   -7.098358E-2   8.381375E-5   1.445279E-6   -1.445279E-6   8.381375E-5   8.382621E-5   9.879071E-1   9.098791E+1   
8.063910E+2   1.100040E+2   1.100040E+2   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   6.485139E-2   -7.161558E-2   8.673663E-5   -1.145863E-6   1.145863E-6   8.673663E-5   8.674420E-5   -7.568806E-1   8.924312E+1   
8.286900E+2   1.099792E+2   1.099792E+2   1.147000E+3   1.147000E+3   9.000000E+1   1.149000E+3   1.149000E+3   6.530699E-2   -7.424999E-2   8.873407E-5   2.394735E-7   -2.394735E-7   8.873407E-5   8.873439E-5   1.546282E-1   9.015463E+1   
8.509110E+2   1.100512E+2   1.100512E+2   1.097000E+3   1.097000E+3   9.000000E+1   1.098000E+3   1.098000E+3   6.543706E-2   -7.572689E-2   8.977637E-5   1.108819E-6   -1.108819E-6   8.977637E-5   8.978322E-5   7.076182E-1   9.070762E+1   
8.732340E+2   1.100229E+2   1.100229E+2   1.047000E+3   1.047000E+3   9.000000E+1   1.048000E+3   1.048000E+3   6.566746E-2   -7.801157E-2   9.140680E-5   2.432068E-6   -2.432068E-6   9.140680E-5   9.143915E-5   1.524114E+0   9.152411E+1   
8.954130E+2   1.100545E+2   1.100545E+2   9.980000E+2   9.980000E+2   9.000000E+1   9.990000E+2   9.990000E+2   6.749747E-2   -7.999315E-2   9.382879E-5   2.374035E-6   -2.374035E-6   9.382879E-5   9.385882E-5   1.449376E+0   9.144938E+1   
9.173480E+2   1.099881E+2   1.099881E+2   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   6.943455E-2   -8.085368E-2   9.558684E-5   1.503901E-6   -1.503901E-6   9.558684E-5   9.559867E-5   9.013803E-1   9.090138E+1   
9.391830E+2   1.100914E+2   1.100914E+2   8.970000E+2   8.970000E+2   9.000000E+1   8.980000E+2   8.980000E+2   7.154162E-2   -8.272604E-2   9.810897E-5   1.169539E-6   -1.169539E-6   9.810897E-5   9.811594E-5   6.829804E-1   9.068298E+1   
9.611110E+2   1.099642E+2   1.099642E+2   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   7.152903E-2   -8.361575E-2   9.868064E-5   1.760521E-6   -1.760521E-6   9.868064E-5   9.869635E-5   1.022082E+0   9.102208E+1   
9.829370E+2   1.100368E+2   1.100368E+2   7.980000E+2   7.980000E+2   9.000000E+1   7.980000E+2   7.980000E+2   7.300593E-2   -8.670946E-2   1.016086E-4   2.690745E-6   -2.690745E-6   1.016086E-4   1.016443E-4   1.516921E+0   9.151692E+1   
1.004828E+3   1.099879E+2   1.099879E+2   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   7.436443E-2   -8.759946E-2   1.030282E-4   2.267812E-6   -2.267812E-6   1.030282E-4   1.030531E-4   1.260966E+0   9.126097E+1   
1.026698E+3   1.100641E+2   1.100641E+2   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   7.500929E-2   -9.002988E-2   1.050098E-4   3.379791E-6   -3.379791E-6   1.050098E-4   1.050641E-4   1.843456E+0   9.184346E+1   
1.048582E+3   1.099921E+2   1.099921E+2   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   7.582014E-2   -9.224069E-2   1.069509E-4   4.225430E-6   -4.225430E-6   1.069509E-4   1.070344E-4   2.262471E+0   9.226247E+1   
1.070415E+3   1.100256E+2   1.100256E+2   5.980000E+2   5.980000E+2   9.000000E+1   5.990000E+2   5.990000E+2   7.741394E-2   -9.310405E-2   1.084986E-4   3.611046E-6   -3.611046E-6   1.084986E-4   1.085587E-4   1.906212E+0   9.190621E+1   
1.092294E+3   1.100245E+2   1.100245E+2   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   7.940441E-2   -9.394625E-2   1.102777E-4   2.689437E-6   -2.689437E-6   1.102777E-4   1.103105E-4   1.397044E+0   9.139704E+1   
1.114129E+3   1.100618E+2   1.100618E+2   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   7.884328E-2   -9.506271E-2   1.106579E-4   3.834378E-6   -3.834378E-6   1.106579E-4   1.107243E-4   1.984546E+0   9.198455E+1   
1.136050E+3   1.100563E+2   1.100563E+2   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   8.152403E-2   -9.772732E-2   1.140507E-4   3.593659E-6   -3.593659E-6   1.140507E-4   1.141073E-4   1.804753E+0   9.180475E+1   
1.157863E+3   1.099824E+2   1.099824E+2   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   8.152926E-2   -9.968804E-2   1.153310E-4   4.871649E-6   -4.871649E-6   1.153310E-4   1.154338E-4   2.418770E+0   9.241877E+1   
1.179952E+3   1.100131E+2   1.100131E+2   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   8.356910E-2   -1.012852E-1   1.176323E-4   4.407105E-6   -4.407105E-6   1.176323E-4   1.177148E-4   2.145588E+0   9.214559E+1   
1.201728E+3   1.100311E+2   1.100311E+2   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   8.345438E-2   -1.023421E-1   1.182497E-4   5.182936E-6   -5.182936E-6   1.182497E-4   1.183633E-4   2.509692E+0   9.250969E+1   
1.223823E+3   1.100265E+2   1.100265E+2   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   8.484996E-2   -1.039856E-1   1.201829E-4   5.225193E-6   -5.225193E-6   1.201829E-4   1.202965E-4   2.489480E+0   9.248948E+1   
1.246112E+3   1.099766E+2   1.099766E+2   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   8.590473E-2   -1.068566E-1   1.227049E-4   6.322006E-6   -6.322006E-6   1.227049E-4   1.228676E-4   2.949388E+0   9.294939E+1   
1.267915E+3   1.099711E+2   1.099711E+2   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   8.746416E-2   -1.076588E-1   1.241915E-4   5.693088E-6   -5.693088E-6   1.241915E-4   1.243219E-4   2.624670E+0   9.262467E+1   
1.289716E+3   1.101041E+2   1.101041E+2   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   8.918069E-2   -1.096873E-1   1.265739E-4   5.749672E-6   -5.749672E-6   1.265739E-4   1.267044E-4   2.600897E+0   9.260090E+1   
1.311406E+3   1.100179E+2   1.100179E+2   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   9.017163E-2   -1.106022E-1   1.277824E-4   5.614847E-6   -5.614847E-6   1.277824E-4   1.279057E-4   2.515999E+0   9.251600E+1   
1.344591E+3   1.101019E+2   1.101019E+2   4.600000E+1   4.600000E+1   9.000000E+1   4.700000E+1   4.700000E+1   8.992344E-2   -1.112103E-1   1.280249E-4   6.195958E-6   -6.195958E-6   1.280249E-4   1.281748E-4   2.770753E+0   9.277075E+1   
1.363608E+3   1.099996E+2   1.099996E+2   4.700000E+1   4.700000E+1   9.000000E+1   4.700000E+1   4.700000E+1   8.867232E-2   -1.110918E-1   1.271743E-4   7.043904E-6   -7.043904E-6   1.271743E-4   1.273692E-4   3.170248E+0   9.317025E+1   
1.385644E+3   1.100554E+2   1.100554E+2   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   8.994245E-2   -1.118321E-1   1.284417E-4   6.588455E-6   -6.588455E-6   1.284417E-4   1.286106E-4   2.936430E+0   9.293643E+1   
1.404692E+3   1.100475E+2   1.100475E+2   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   9.036919E-2   -1.120162E-1   1.288254E-4   6.393180E-6   -6.393180E-6   1.288254E-4   1.289840E-4   2.841069E+0   9.284107E+1   
1.427118E+3   1.099919E+2   1.099919E+2   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   9.026551E-2   -1.110059E-1   1.281033E-4   5.809371E-6   -5.809371E-6   1.281033E-4   1.282350E-4   2.596533E+0   9.259653E+1   
1.446186E+3   1.099965E+2   1.099965E+2   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   8.962183E-2   -1.110611E-1   1.277414E-4   6.321546E-6   -6.321546E-6   1.277414E-4   1.278977E-4   2.833089E+0   9.283309E+1   
1.468542E+3   1.099915E+2   1.099915E+2   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   9.054529E-2   -1.112790E-1   1.284542E-4   5.780949E-6   -5.780949E-6   1.284542E-4   1.285842E-4   2.576800E+0   9.257680E+1   
1.487625E+3   1.099992E+2   1.099992E+2   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   8.948439E-2   -1.115800E-1   1.279943E-4   6.762389E-6   -6.762389E-6   1.279943E-4   1.281728E-4   3.024326E+0   9.302433E+1   
1.510059E+3   1.100657E+2   1.100657E+2   3.100000E+1   3.100000E+1   9.000000E+1   3.100000E+1   3.100000E+1   9.081961E-2   -1.112692E-1   1.286174E-4   5.571648E-6   -5.571648E-6   1.286174E-4   1.287380E-4   2.480477E+0   9.248048E+1   
1.531480E+3   1.100645E+2   1.100645E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   8.905028E-2   -1.113873E-1   1.276004E-4   6.957494E-6   -6.957494E-6   1.276004E-4   1.277899E-4   3.120999E+0   9.312100E+1   
1.550544E+3   1.100088E+2   1.100088E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   9.061709E-2   -1.127574E-1   1.294614E-4   6.694406E-6   -6.694406E-6   1.294614E-4   1.296344E-4   2.960108E+0   9.296011E+1   
1.572974E+3   1.099875E+2   1.099875E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   9.155343E-2   -1.108025E-1   1.287671E-4   4.723811E-6   -4.723811E-6   1.287671E-4   1.288537E-4   2.100948E+0   9.210095E+1   
1.592007E+3   1.100121E+2   1.100121E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   8.977433E-2   -1.122494E-1   1.286095E-4   6.985584E-6   -6.985584E-6   1.286095E-4   1.287991E-4   3.109036E+0   9.310904E+1   
1.614455E+3   1.099967E+2   1.099967E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   9.034987E-2   -1.121687E-1   1.289128E-4   6.507142E-6   -6.507142E-6   1.289128E-4   1.290769E-4   2.889671E+0   9.288967E+1   
1.633499E+3   1.100055E+2   1.100055E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   9.107667E-2   -1.111799E-1   1.287181E-4   5.323131E-6   -5.323131E-6   1.287181E-4   1.288282E-4   2.368114E+0   9.236811E+1   
1.655967E+3   1.099988E+2   1.099988E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   9.060729E-2   -1.120030E-1   1.289640E-4   6.208439E-6   -6.208439E-6   1.289640E-4   1.291134E-4   2.756140E+0   9.275614E+1   
1.674989E+3   1.100189E+2   1.100189E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   9.142334E-2   -1.113216E-1   1.290248E-4   5.159389E-6   -5.159389E-6   1.290248E-4   1.291279E-4   2.289900E+0   9.228990E+1   
1.697401E+3   1.099978E+2   1.099978E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   9.227379E-2   -1.123077E-1   1.301928E-4   5.175018E-6   -5.175018E-6   1.301928E-4   1.302956E-4   2.276245E+0   9.227625E+1   
1.716463E+3   1.100551E+2   1.100551E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   9.155071E-2   -1.122632E-1   1.297167E-4   5.680742E-6   -5.680742E-6   1.297167E-4   1.298411E-4   2.507577E+0   9.250758E+1   
1.738567E+3   1.100205E+2   1.100205E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   9.154852E-2   -1.121616E-1   1.296493E-4   5.615972E-6   -5.615972E-6   1.296493E-4   1.297708E-4   2.480311E+0   9.248031E+1   
1.757235E+3   1.100460E+2   1.100460E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   9.130400E-2   -1.121758E-1   1.295073E-4   5.806063E-6   -5.806063E-6   1.295073E-4   1.296374E-4   2.566962E+0   9.256696E+1   
1.779212E+3   1.099858E+2   1.099858E+2   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   9.056890E-2   -1.132176E-1   1.297314E-4   7.030897E-6   -7.030897E-6   1.297314E-4   1.299217E-4   3.102157E+0   9.310216E+1   
1.797889E+3   1.100472E+2   1.100472E+2   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   9.156910E-2   -1.115815E-1   1.292841E-4   5.221479E-6   -5.221479E-6   1.292841E-4   1.293895E-4   2.312783E+0   9.231278E+1   
1.819901E+3   1.099804E+2   1.099804E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   9.201763E-2   -1.125924E-1   1.302198E-4   5.550612E-6   -5.550612E-6   1.302198E-4   1.303381E-4   2.440752E+0   9.244075E+1   
1.838614E+3   1.099953E+2   1.099953E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   9.086467E-2   -1.127783E-1   1.296281E-4   6.524925E-6   -6.524925E-6   1.296281E-4   1.297922E-4   2.881593E+0   9.288159E+1   
1.860674E+3   1.100019E+2   1.100019E+2   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   9.159547E-2   -1.132185E-1   1.303666E-4   6.272207E-6   -6.272207E-6   1.303666E-4   1.305174E-4   2.754494E+0   9.275449E+1   
1.882701E+3   1.099852E+2   1.099852E+2   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   9.063674E-2   -1.132719E-1   1.298087E-4   7.016223E-6   -7.016223E-6   1.298087E-4   1.299981E-4   3.093855E+0   9.309386E+1   
1.904779E+3   1.099654E+2   1.099654E+2   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   9.045547E-2   -1.130483E-1   1.295509E-4   7.004085E-6   -7.004085E-6   1.295509E-4   1.297401E-4   3.094645E+0   9.309465E+1   
1.926906E+3   1.100355E+2   1.100355E+2   -8.000000E+0   -8.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   9.150893E-2   -1.134777E-1   1.304820E-4   6.505697E-6   -6.505697E-6   1.304820E-4   1.306440E-4   2.854346E+0   9.285435E+1   
1.949039E+3   1.099769E+2   1.099769E+2   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   9.066065E-2   -1.141141E-1   1.303719E-4   7.549119E-6   -7.549119E-6   1.303719E-4   1.305903E-4   3.313982E+0   9.331398E+1   
1.971216E+3   1.099993E+2   1.099993E+2   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   9.127672E-2   -1.144751E-1   1.309880E-4   7.329525E-6   -7.329525E-6   1.309880E-4   1.311929E-4   3.202686E+0   9.320269E+1   
1.993499E+3   1.100576E+2   1.100576E+2   -1.300000E+1   -1.300000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   9.199092E-2   -1.131949E-1   1.305957E-4   5.964291E-6   -5.964291E-6   1.305957E-4   1.307319E-4   2.614874E+0   9.261487E+1   
2.015431E+3   1.099659E+2   1.099659E+2   -1.500000E+1   -1.500000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   9.201520E-2   -1.131621E-1   1.305894E-4   5.924869E-6   -5.924869E-6   1.305894E-4   1.307237E-4   2.597741E+0   9.259774E+1   
2.037286E+3   1.099859E+2   1.099859E+2   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   9.172926E-2   -1.129952E-1   1.303039E-4   6.027245E-6   -6.027245E-6   1.303039E-4   1.304432E-4   2.648346E+0   9.264835E+1   
2.059478E+3   1.099956E+2   1.099956E+2   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   9.246587E-2   -1.135339E-1   1.311102E-4   5.834643E-6   -5.834643E-6   1.311102E-4   1.312399E-4   2.548086E+0   9.254809E+1   
2.081751E+3   1.100607E+2   1.100607E+2   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   9.160930E-2   -1.137290E-1   1.307077E-4   6.595753E-6   -6.595753E-6   1.307077E-4   1.308740E-4   2.888801E+0   9.288880E+1   
2.104037E+3   1.100564E+2   1.100564E+2   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.200000E+1   -2.200000E+1   9.093739E-2   -1.135186E-1   1.301552E-4   6.955131E-6   -6.955131E-6   1.301552E-4   1.303409E-4   3.058818E+0   9.305882E+1   
2.126237E+3   1.100354E+2   1.100354E+2   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   9.341483E-2   -1.137088E-1   1.318107E-4   5.247085E-6   -5.247085E-6   1.318107E-4   1.319151E-4   2.279610E+0   9.227961E+1   
2.148528E+3   1.100192E+2   1.100192E+2   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   9.221186E-2   -1.129498E-1   1.305727E-4   5.640624E-6   -5.640624E-6   1.305727E-4   1.306945E-4   2.473589E+0   9.247359E+1   
2.170753E+3   1.100450E+2   1.100450E+2   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   9.174153E-2   -1.134189E-1   1.305874E-4   6.295165E-6   -6.295165E-6   1.305874E-4   1.307391E-4   2.759894E+0   9.275989E+1   
2.193026E+3   1.099948E+2   1.099948E+2   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   9.102606E-2   -1.137701E-1   1.303738E-4   7.053996E-6   -7.053996E-6   1.303738E-4   1.305645E-4   3.097020E+0   9.309702E+1   
2.215305E+3   1.100064E+2   1.100064E+2   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   9.222969E-2   -1.145764E-1   1.316431E-4   6.690862E-6   -6.690862E-6   1.316431E-4   1.318130E-4   2.909599E+0   9.290960E+1   
2.237576E+3   1.100006E+2   1.100006E+2   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   9.273863E-2   -1.146012E-1   1.319739E-4   6.330682E-6   -6.330682E-6   1.319739E-4   1.321257E-4   2.746327E+0   9.274633E+1   
2.259847E+3   1.100128E+2   1.100128E+2   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   9.204529E-2   -1.141128E-1   1.312272E-4   6.524190E-6   -6.524190E-6   1.312272E-4   1.313893E-4   2.846217E+0   9.284622E+1   
2.282126E+3   1.100294E+2   1.100294E+2   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   9.207102E-2   -1.145574E-1   1.315326E-4   6.795787E-6   -6.795787E-6   1.315326E-4   1.317080E-4   2.957624E+0   9.295762E+1   
2.304370E+3   1.100404E+2   1.100404E+2   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   9.255452E-2   -1.143475E-1   1.316949E-4   6.300987E-6   -6.300987E-6   1.316949E-4   1.318455E-4   2.739248E+0   9.273925E+1   
2.326650E+3   1.100200E+2   1.100200E+2   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   9.294790E-2   -1.147273E-1   1.321854E-4   6.258332E-6   -6.258332E-6   1.321854E-4   1.323335E-4   2.710650E+0   9.271065E+1   
2.348903E+3   1.100246E+2   1.100246E+2   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   9.119110E-2   -1.133290E-1   1.301886E-4   6.643510E-6   -6.643510E-6   1.301886E-4   1.303580E-4   2.921264E+0   9.292126E+1   
2.371127E+3   1.100498E+2   1.100498E+2   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   9.230205E-2   -1.150657E-1   1.320065E-4   6.957254E-6   -6.957254E-6   1.320065E-4   1.321897E-4   3.016917E+0   9.301692E+1   
2.393363E+3   1.099953E+2   1.099953E+2   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   9.172250E-2   -1.135321E-1   1.306494E-4   6.383250E-6   -6.383250E-6   1.306494E-4   1.308052E-4   2.797125E+0   9.279713E+1   
2.426695E+3   1.100470E+2   1.100470E+2   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   9.197348E-2   -1.173182E-1   1.332704E-4   8.672878E-6   -8.672878E-6   1.332704E-4   1.335523E-4   3.723404E+0   9.372340E+1   
2.448414E+3   1.099721E+2   1.099721E+2   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   9.423648E-2   -1.173802E-1   1.347099E-4   7.039619E-6   -7.039619E-6   1.347099E-4   1.348937E-4   2.991421E+0   9.299142E+1   
2.470154E+3   1.100021E+2   1.100021E+2   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   9.639731E-2   -1.197621E-1   1.375971E-4   6.998636E-6   -6.998636E-6   1.375971E-4   1.377750E-4   2.911740E+0   9.291174E+1   
2.491914E+3   1.100317E+2   1.100317E+2   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   9.744936E-2   -1.198198E-1   1.382851E-4   6.258211E-6   -6.258211E-6   1.382851E-4   1.384266E-4   2.591202E+0   9.259120E+1   
2.514093E+3   1.100332E+2   1.100332E+2   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   9.832369E-2   -1.217532E-1   1.400849E-4   6.875536E-6   -6.875536E-6   1.400849E-4   1.402535E-4   2.809892E+0   9.280989E+1   
2.535767E+3   1.099347E+2   1.099347E+2   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   9.846054E-2   -1.239731E-1   1.416153E-4   8.225657E-6   -8.225657E-6   1.416153E-4   1.418540E-4   3.324263E+0   9.332426E+1   
2.557504E+3   1.100883E+2   1.100883E+2   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   9.938157E-2   -1.256516E-1   1.432779E-4   8.641757E-6   -8.641757E-6   1.432779E-4   1.435383E-4   3.451594E+0   9.345159E+1   
2.579941E+3   1.099988E+2   1.099988E+2   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   1.010889E-1   -1.254641E-1   1.442113E-4   7.256448E-6   -7.256448E-6   1.442113E-4   1.443938E-4   2.880588E+0   9.288059E+1   
2.601638E+3   1.100344E+2   1.100344E+2   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   1.018816E-1   -1.285539E-1   1.467137E-4   8.690080E-6   -8.690080E-6   1.467137E-4   1.469709E-4   3.389757E+0   9.338976E+1   
2.623299E+3   1.100048E+2   1.100048E+2   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   1.018620E-1   -1.296838E-1   1.474375E-4   9.443299E-6   -9.443299E-6   1.474375E-4   1.477396E-4   3.664760E+0   9.366476E+1   
2.644997E+3   1.100341E+2   1.100341E+2   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   1.038663E-1   -1.309027E-1   1.494705E-4   8.757744E-6   -8.757744E-6   1.494705E-4   1.497268E-4   3.353229E+0   9.335323E+1   
2.666722E+3   1.100461E+2   1.100461E+2   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.500000E+2   -6.500000E+2   1.041071E-1   -1.323587E-1   1.505677E-4   9.531541E-6   -9.531541E-6   1.505677E-4   1.508691E-4   3.622220E+0   9.362222E+1   
2.688352E+3   1.099203E+2   1.099203E+2   -7.000000E+2   -7.000000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   1.046154E-1   -1.347689E-1   1.524517E-4   1.073124E-5   -1.073124E-5   1.524517E-4   1.528289E-4   4.026469E+0   9.402647E+1   
2.710075E+3   1.099821E+2   1.099821E+2   -7.500000E+2   -7.500000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   1.056613E-1   -1.363728E-1   1.541429E-4   1.100629E-5   -1.100629E-5   1.541429E-4   1.545353E-4   4.084169E+0   9.408417E+1   
2.731710E+3   1.100285E+2   1.100285E+2   -8.000000E+2   -8.000000E+2   9.000000E+1   -8.000000E+2   -8.000000E+2   1.069428E-1   -1.368290E-1   1.552323E-4   1.035673E-5   -1.035673E-5   1.552323E-4   1.555774E-4   3.816981E+0   9.381698E+1   
2.753425E+3   1.099886E+2   1.099886E+2   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   1.070336E-1   -1.393385E-1   1.569229E-4   1.193025E-5   -1.193025E-5   1.569229E-4   1.573757E-4   4.347617E+0   9.434762E+1   
2.775141E+3   1.099837E+2   1.099837E+2   -9.000000E+2   -9.000000E+2   9.000000E+1   -8.990000E+2   -8.990000E+2   1.106688E-1   -1.401540E-1   1.597014E-4   9.774667E-6   -9.774667E-6   1.597014E-4   1.600003E-4   3.502470E+0   9.350247E+1   
2.796869E+3   1.100590E+2   1.100590E+2   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.490000E+2   -9.490000E+2   1.105721E-1   -1.407387E-1   1.600225E-4   1.022842E-5   -1.022842E-5   1.600225E-4   1.603491E-4   3.657292E+0   9.365729E+1   
2.818604E+3   1.100328E+2   1.100328E+2   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   1.120727E-1   -1.435155E-1   1.627587E-4   1.093396E-5   -1.093396E-5   1.627587E-4   1.631255E-4   3.843297E+0   9.384330E+1   
2.840732E+3   1.100352E+2   1.100352E+2   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   1.128040E-1   -1.441819E-1   1.636449E-4   1.082865E-5   -1.082865E-5   1.636449E-4   1.640027E-4   3.785839E+0   9.378584E+1   
2.862504E+3   1.100413E+2   1.100413E+2   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   1.142770E-1   -1.453526E-1   1.653180E-4   1.050462E-5   -1.050462E-5   1.653180E-4   1.656514E-4   3.635796E+0   9.363580E+1   
2.884367E+3   1.099746E+2   1.099746E+2   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.150000E+3   -1.150000E+3   1.133072E-1   -1.486273E-1   1.668512E-4   1.336281E-5   -1.336281E-5   1.668512E-4   1.673854E-4   4.578943E+0   9.457894E+1   
2.906945E+3   1.100378E+2   1.100378E+2   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   1.156066E-1   -1.485917E-1   1.682496E-4   1.163883E-5   -1.163883E-5   1.682496E-4   1.686517E-4   3.957185E+0   9.395719E+1   
2.928785E+3   1.099757E+2   1.099757E+2   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   1.149249E-1   -1.508730E-1   1.693139E-4   1.363450E-5   -1.363450E-5   1.693139E-4   1.698620E-4   4.603974E+0   9.460397E+1   
2.950659E+3   1.100229E+2   1.100229E+2   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   1.176409E-1   -1.518830E-1   1.716509E-4   1.228591E-5   -1.228591E-5   1.716509E-4   1.720900E-4   4.093962E+0   9.409396E+1   
2.973281E+3   1.100366E+2   1.100366E+2   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   1.189976E-1   -1.540428E-1   1.738963E-4   1.269453E-5   -1.269453E-5   1.738963E-4   1.743590E-4   4.175218E+0   9.417522E+1   
2.995122E+3   1.100582E+2   1.100582E+2   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   1.181008E-1   -1.558876E-1   1.745434E-4   1.456384E-5   -1.456384E-5   1.745434E-4   1.751499E-4   4.769692E+0   9.476969E+1   
3.016992E+3   1.099996E+2   1.099996E+2   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   1.208742E-1   -1.567653E-1   1.768297E-4   1.308638E-5   -1.308638E-5   1.768297E-4   1.773132E-4   4.232492E+0   9.423249E+1   
3.039397E+3   1.099294E+2   1.099294E+2   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   1.213050E-1   -1.594770E-1   1.788621E-4   1.454065E-5   -1.454065E-5   1.788621E-4   1.794522E-4   4.647656E+0   9.464766E+1   
3.061250E+3   1.100014E+2   1.100014E+2   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.548000E+3   -1.548000E+3   1.224343E-1   -1.610174E-1   1.805635E-4   1.471245E-5   -1.471245E-5   1.805635E-4   1.811619E-4   4.658213E+0   9.465821E+1   
3.083385E+3   1.099936E+2   1.099936E+2   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   1.232482E-1   -1.624603E-1   1.820064E-4   1.505375E-5   -1.505375E-5   1.820064E-4   1.826279E-4   4.728170E+0   9.472817E+1   
3.106260E+3   1.100222E+2   1.100222E+2   -1.650000E+3   -1.650000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   1.250147E-1   -1.640261E-1   1.841184E-4   1.477090E-5   -1.477090E-5   1.841184E-4   1.847100E-4   4.586731E+0   9.458673E+1   
3.128305E+3   1.100712E+2   1.100712E+2   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.698000E+3   -1.698000E+3   1.252850E-1   -1.652613E-1   1.850900E-4   1.537849E-5   -1.537849E-5   1.850900E-4   1.857277E-4   4.749599E+0   9.474960E+1   
3.150453E+3   1.099966E+2   1.099966E+2   -1.750000E+3   -1.750000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   1.260655E-1   -1.678887E-1   1.872837E-4   1.651891E-5   -1.651891E-5   1.872837E-4   1.880108E-4   5.040594E+0   9.504059E+1   
3.173646E+3   1.100724E+2   1.100724E+2   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.798000E+3   -1.798000E+3   1.270187E-1   -1.680049E-1   1.879487E-4   1.588992E-5   -1.588992E-5   1.879487E-4   1.886192E-4   4.832518E+0   9.483252E+1   
3.195785E+3   1.099422E+2   1.099422E+2   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.848000E+3   -1.848000E+3   1.284023E-1   -1.706038E-1   1.904967E-4   1.656559E-5   -1.656559E-5   1.904967E-4   1.912157E-4   4.969937E+0   9.496994E+1   
3.217911E+3   1.100013E+2   1.100013E+2   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   1.288732E-1   -1.703445E-1   1.906190E-4   1.604780E-5   -1.604780E-5   1.906190E-4   1.912934E-4   4.812258E+0   9.481226E+1   
3.241070E+3   1.100113E+2   1.100113E+2   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.948000E+3   -1.948000E+3   1.297810E-1   -1.729741E-1   1.928929E-4   1.709548E-5   -1.709548E-5   1.928929E-4   1.936490E-4   5.064708E+0   9.506471E+1   
3.263558E+3   1.100119E+2   1.100119E+2   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   1.303787E-1   -1.748326E-1   1.944728E-4   1.786850E-5   -1.786850E-5   1.944728E-4   1.952920E-4   5.249697E+0   9.524970E+1   
3.301058E+3   1.100387E+2   1.100387E+2   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.415950E-1   -1.920734E-1   2.126360E-4   2.084411E-5   -2.084411E-5   2.126360E-4   2.136552E-4   5.598657E+0   9.559866E+1   
3.327165E+3   1.099546E+2   1.099546E+2   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.500398E-1   -2.093079E-1   2.290816E-4   2.586550E-5   -2.586550E-5   2.290816E-4   2.305372E-4   6.441958E+0   9.644196E+1   
3.352348E+3   1.100585E+2   1.100585E+2   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.616006E-1   -2.253455E-1   2.466742E-4   2.779965E-5   -2.779965E-5   2.466742E-4   2.482357E-4   6.429980E+0   9.642998E+1   
3.378041E+3   1.100884E+2   1.100884E+2   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   1.720500E-1   -2.395699E-1   2.623987E-4   2.937053E-5   -2.937053E-5   2.623987E-4   2.640373E-4   6.386587E+0   9.638659E+1   
3.403809E+3   1.100639E+2   1.100639E+2   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   1.764224E-1   -2.504727E-1   2.722028E-4   3.326448E-5   -3.326448E-5   2.722028E-4   2.742278E-4   6.967273E+0   9.696727E+1   
3.428534E+3   1.099770E+2   1.099770E+2   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   1.761524E-1   -2.527528E-1   2.735209E-4   3.495483E-5   -3.495483E-5   2.735209E-4   2.757454E-4   7.282688E+0   9.728269E+1   
3.453780E+3   1.100683E+2   1.100683E+2   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   1.646170E-1   -2.400108E-1   2.580904E-4   3.515643E-5   -3.515643E-5   2.580904E-4   2.604739E-4   7.756945E+0   9.775694E+1   
3.479467E+3   1.100019E+2   1.100019E+2   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   1.448525E-1   -2.217075E-1   2.339504E-4   3.780869E-5   -3.780869E-5   2.339504E-4   2.369858E-4   9.180190E+0   9.918019E+1   
3.504200E+3   1.099878E+2   1.099878E+2   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.299645E-1   -2.056061E-1   2.142592E-4   3.829372E-5   -3.829372E-5   2.142592E-4   2.176544E-4   1.013326E+1   1.001333E+2   
3.528847E+3   1.100875E+2   1.100875E+2   -7.000000E+3   -7.000000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.222769E-1   -1.976593E-1   2.043307E-4   3.878428E-5   -3.878428E-5   2.043307E-4   2.079790E-4   1.074753E+1   1.007475E+2   
3.554045E+3   1.100571E+2   1.100571E+2   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.183466E-1   -1.944971E-1   1.998413E-4   3.962392E-5   -3.962392E-5   1.998413E-4   2.037317E-4   1.121497E+1   1.012150E+2   
3.579243E+3   1.100456E+2   1.100456E+2   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.245616E-1   -2.015172E-1   2.082558E-4   3.961665E-5   -3.961665E-5   2.082558E-4   2.119905E-4   1.077072E+1   1.007707E+2   
3.604444E+3   1.099893E+2   1.099893E+2   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.325149E-1   -2.147357E-1   2.217819E-4   4.237601E-5   -4.237601E-5   2.217819E-4   2.257941E-4   1.081716E+1   1.008172E+2   
3.630044E+3   1.100122E+2   1.100122E+2   -9.000000E+3   -9.000000E+3   9.000000E+1   -9.000000E+3   -9.000000E+3   1.453922E-1   -2.319679E-1   2.409665E-4   4.411748E-5   -4.411748E-5   2.409665E-4   2.449718E-4   1.037512E+1   1.003751E+2   
3.655248E+3   1.099813E+2   1.099813E+2   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.553991E-1   -2.506426E-1   2.593159E-4   4.892504E-5   -4.892504E-5   2.593159E-4   2.638909E-4   1.068438E+1   1.006844E+2   
3.680482E+3   1.099977E+2   1.099977E+2   -9.999000E+3   -9.999000E+3   9.000000E+1   -9.998000E+3   -9.998000E+3   1.654220E-1   -2.634333E-1   2.738429E-4   4.987396E-5   -4.987396E-5   2.738429E-4   2.783476E-4   1.032193E+1   1.003219E+2   
3.717071E+3   1.099942E+2   1.099942E+2   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.419635E-1   -2.345315E-1   2.405163E-4   4.832945E-5   -4.832945E-5   2.405163E-4   2.453239E-4   1.136173E+1   1.013617E+2   
3.741666E+3   1.099922E+2   1.099922E+2   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.282860E-1   -2.156981E-1   2.197943E-4   4.613299E-5   -4.613299E-5   2.197943E-4   2.245836E-4   1.185383E+1   1.018538E+2   
3.765919E+3   1.100405E+2   1.100405E+2   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.137468E-1   -1.976697E-1   1.990638E-4   4.510019E-5   -4.510019E-5   1.990638E-4   2.041088E-4   1.276551E+1   1.027655E+2   
3.790569E+3   1.100649E+2   1.100649E+2   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.026817E-1   -1.788301E-1   1.799528E-4   4.096748E-5   -4.096748E-5   1.799528E-4   1.845572E-4   1.282519E+1   1.028252E+2   
3.815273E+3   1.100077E+2   1.100077E+2   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   8.854014E-2   -1.618123E-1   1.601263E-4   4.030128E-5   -4.030128E-5   1.601263E-4   1.651200E-4   1.412704E+1   1.041270E+2   
3.840473E+3   1.100281E+2   1.100281E+2   -7.000000E+3   -7.000000E+3   9.000000E+1   -6.999000E+3   -6.999000E+3   8.137738E-2   -1.454504E-1   1.450416E-4   3.490216E-5   -3.490216E-5   1.450416E-4   1.491819E-4   1.353015E+1   1.035302E+2   
3.865164E+3   1.100000E+2   1.100000E+2   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   6.796225E-2   -1.267944E-1   1.245973E-4   3.262760E-5   -3.262760E-5   1.245973E-4   1.287985E-4   1.467423E+1   1.046742E+2   
3.889354E+3   1.100420E+2   1.100420E+2   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   5.798843E-2   -1.105028E-1   1.078205E-4   2.935355E-5   -2.935355E-5   1.078205E-4   1.117447E-4   1.522938E+1   1.052294E+2   
3.914061E+3   1.099981E+2   1.099981E+2   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   4.509752E-2   -9.223672E-2   8.795420E-5   2.694624E-5   -2.694624E-5   8.795420E-5   9.198935E-5   1.703332E+1   1.070333E+2   
3.939216E+3   1.100110E+2   1.100110E+2   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   3.672601E-2   -7.723723E-2   7.300952E-5   2.333182E-5   -2.333182E-5   7.300952E-5   7.664701E-5   1.772244E+1   1.077224E+2   
3.963908E+3   1.099962E+2   1.099962E+2   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   2.491018E-2   -5.973809E-2   5.430742E-5   2.063074E-5   -2.063074E-5   5.430742E-5   5.809409E-5   2.080118E+1   1.108012E+2   
3.988598E+3   1.100669E+2   1.100669E+2   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   1.425918E-2   -4.218600E-2   3.629099E-5   1.703348E-5   -1.703348E-5   3.629099E-5   4.008959E-5   2.514341E+1   1.151434E+2   
4.013302E+3   1.099981E+2   1.099981E+2   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   2.847970E-3   -2.742313E-2   1.962114E-5   1.582202E-5   -1.582202E-5   1.962114E-5   2.520566E-5   3.888188E+1   1.288819E+2   
4.037501E+3   1.100680E+2   1.100680E+2   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   -8.954403E-3   -8.360448E-3   -9.096025E-8   1.208878E-5   -1.208878E-5   -9.096025E-8   1.208912E-5   9.043111E+1   1.804311E+2   
4.062704E+3   1.100127E+2   1.100127E+2   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   -1.824106E-2   7.395274E-3   -1.609394E-5   8.656834E-6   -8.656834E-6   -1.609394E-5   1.827446E-5   1.517245E+2   2.417245E+2   
4.087409E+3   1.100241E+2   1.100241E+2   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   -3.075582E-2   2.505990E-2   -3.533593E-5   6.364505E-6   -6.364505E-6   -3.533593E-5   3.590453E-5   1.697897E+2   2.597897E+2   
4.121066E+3   1.100967E+2   1.100967E+2   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   -3.026435E-2   2.749769E-2   -3.661979E-5   4.407242E-6   -4.407242E-6   -3.661979E-5   3.688405E-5   1.731374E+2   2.631374E+2   
4.143061E+3   1.100166E+2   1.100166E+2   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.899000E+3   -1.899000E+3   -3.093438E-2   2.963849E-2   -3.842832E-5   3.503221E-6   -3.503221E-6   -3.842832E-5   3.858767E-5   1.747912E+2   2.647912E+2   
4.165108E+3   1.099805E+2   1.099805E+2   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.849000E+3   -1.849000E+3   -3.198115E-2   3.127093E-2   -4.013867E-5   3.210205E-6   -3.210205E-6   -4.013867E-5   4.026684E-5   1.754273E+2   2.654273E+2   
4.186894E+3   1.099586E+2   1.099586E+2   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.799000E+3   -1.799000E+3   -3.250607E-2   3.272850E-2   -4.141250E-5   2.645528E-6   -2.645528E-6   -4.141250E-5   4.149692E-5   1.763448E+2   2.663448E+2   
4.208931E+3   1.099892E+2   1.099892E+2   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   -3.488801E-2   3.520770E-2   -4.449980E-5   2.786455E-6   -2.786455E-6   -4.449980E-5   4.458695E-5   1.764170E+2   2.664170E+2   
4.230955E+3   1.100757E+2   1.100757E+2   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   -3.575777E-2   3.659839E-2   -4.594327E-5   2.520566E-6   -2.520566E-6   -4.594327E-5   4.601236E-5   1.768598E+2   2.668598E+2   
4.252997E+3   1.100423E+2   1.100423E+2   -1.650000E+3   -1.650000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   -3.706900E-2   3.773044E-2   -4.749122E-5   2.750292E-6   -2.750292E-6   -4.749122E-5   4.757079E-5   1.766856E+2   2.666856E+2   
4.274830E+3   1.100009E+2   1.100009E+2   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.599000E+3   -1.599000E+3   -3.722822E-2   3.863028E-2   -4.817572E-5   2.279765E-6   -2.279765E-6   -4.817572E-5   4.822963E-5   1.772907E+2   2.672907E+2   
4.296970E+3   1.100141E+2   1.100141E+2   -1.550000E+3   -1.550000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   -3.862045E-2   3.981479E-2   -4.980792E-5   2.535102E-6   -2.535102E-6   -4.980792E-5   4.987239E-5   1.770863E+2   2.670863E+2   
4.318704E+3   1.100109E+2   1.100109E+2   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   -3.929235E-2   4.369359E-2   -5.274954E-5   4.962045E-7   -4.962045E-7   -5.274954E-5   5.275188E-5   1.794610E+2   2.694610E+2   
4.340829E+3   1.100264E+2   1.100264E+2   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   -4.029094E-2   4.405192E-2   -5.360030E-5   1.000531E-6   -1.000531E-6   -5.360030E-5   5.360963E-5   1.789306E+2   2.689306E+2   
4.362928E+3   1.100547E+2   1.100547E+2   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   -4.136564E-2   4.572704E-2   -5.535571E-5   7.002665E-7   -7.002665E-7   -5.535571E-5   5.536014E-5   1.792752E+2   2.692752E+2   
4.385004E+3   1.099715E+2   1.099715E+2   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   -4.194794E-2   4.725584E-2   -5.671141E-5   1.314666E-7   -1.314666E-7   -5.671141E-5   5.671156E-5   1.798672E+2   2.698672E+2   
4.407127E+3   1.099755E+2   1.099755E+2   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   -4.374760E-2   4.929394E-2   -5.915144E-5   1.301025E-7   -1.301025E-7   -5.915144E-5   5.915158E-5   1.798740E+2   2.698740E+2   
4.429201E+3   1.100178E+2   1.100178E+2   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.250000E+3   -1.250000E+3   -4.450264E-2   5.120893E-2   -6.086544E-5   -5.634176E-7   5.634176E-7   -6.086544E-5   6.086805E-5   -1.794696E+2   -8.946964E+1   
4.451042E+3   1.100177E+2   1.100177E+2   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   -4.452748E-2   5.257447E-2   -6.177016E-5   -1.437794E-6   1.437794E-6   -6.177016E-5   6.178690E-5   -1.786666E+2   -8.866659E+1   
4.473130E+3   1.100257E+2   1.100257E+2   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   -4.533466E-2   5.454654E-2   -6.355359E-5   -2.130063E-6   2.130063E-6   -6.355359E-5   6.358928E-5   -1.780804E+2   -8.808039E+1   
4.495244E+3   1.099995E+2   1.099995E+2   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   -4.617959E-2   5.566142E-2   -6.480208E-5   -2.234001E-6   2.234001E-6   -6.480208E-5   6.484057E-5   -1.780256E+2   -8.802555E+1   
4.517309E+3   1.100428E+2   1.100428E+2   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   -4.820019E-2   5.653392E-2   -6.661956E-5   -1.309920E-6   1.309920E-6   -6.661956E-5   6.663243E-5   -1.788736E+2   -8.887356E+1   
4.539386E+3   1.099523E+2   1.099523E+2   -1.000000E+3   -1.000000E+3   9.000000E+1   -1.000000E+3   -1.000000E+3   -4.859593E-2   5.966844E-2   -6.890570E-5   -3.066480E-6   3.066480E-6   -6.890570E-5   6.897390E-5   -1.774519E+2   -8.745187E+1   
4.561301E+3   1.100138E+2   1.100138E+2   -9.510000E+2   -9.510000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   -4.902821E-2   5.977858E-2   -6.924469E-5   -2.818764E-6   2.818764E-6   -6.924469E-5   6.930203E-5   -1.776689E+2   -8.766893E+1   
4.582984E+3   1.099868E+2   1.099868E+2   -9.000000E+2   -9.000000E+2   9.000000E+1   -9.000000E+2   -9.000000E+2   -5.177771E-2   6.339107E-2   -7.329733E-5   -3.146893E-6   3.146893E-6   -7.329733E-5   7.336486E-5   -1.775416E+2   -8.754162E+1   
4.604842E+3   1.099913E+2   1.099913E+2   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   -5.074752E-2   6.266887E-2   -7.219006E-5   -3.436691E-6   3.436691E-6   -7.219006E-5   7.227182E-5   -1.772744E+2   -8.727443E+1   
4.626469E+3   1.099671E+2   1.099671E+2   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   -5.267696E-2   6.498270E-2   -7.488990E-5   -3.522338E-6   3.522338E-6   -7.488990E-5   7.497269E-5   -1.773072E+2   -8.730716E+1   
4.648193E+3   1.099726E+2   1.099726E+2   -7.510000E+2   -7.510000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   -5.507974E-2   6.492502E-2   -7.633785E-5   -1.707457E-6   1.707457E-6   -7.633785E-5   7.635694E-5   -1.787187E+2   -8.871867E+1   
4.670062E+3   1.100032E+2   1.100032E+2   -7.000000E+2   -7.000000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   -5.516595E-2   6.673203E-2   -7.756803E-5   -2.825065E-6   2.825065E-6   -7.756803E-5   7.761946E-5   -1.779142E+2   -8.791418E+1   
4.692019E+3   1.099926E+2   1.099926E+2   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.490000E+2   -6.490000E+2   -5.547429E-2   6.934160E-2   -7.945825E-5   -4.303069E-6   4.303069E-6   -7.945825E-5   7.957468E-5   -1.769002E+2   -8.690017E+1   
4.713655E+3   1.100132E+2   1.100132E+2   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   -5.794580E-2   7.087189E-2   -8.198292E-5   -3.475525E-6   3.475525E-6   -8.198292E-5   8.205655E-5   -1.775725E+2   -8.757250E+1   
4.735326E+3   1.100177E+2   1.100177E+2   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   -5.750985E-2   7.255618E-2   -8.281035E-5   -4.899107E-6   4.899107E-6   -8.281035E-5   8.295514E-5   -1.766143E+2   -8.661430E+1   
4.757270E+3   1.099909E+2   1.099909E+2   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   -5.912636E-2   7.322252E-2   -8.424373E-5   -4.139124E-6   4.139124E-6   -8.424373E-5   8.434536E-5   -1.771872E+2   -8.718716E+1   
4.778900E+3   1.100002E+2   1.100002E+2   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   -5.942885E-2   7.454112E-2   -8.528954E-5   -4.777456E-6   4.777456E-6   -8.528954E-5   8.542324E-5   -1.767940E+2   -8.679395E+1   
4.800523E+3   1.100012E+2   1.100012E+2   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   -6.045813E-2   7.763820E-2   -8.794298E-5   -6.040950E-6   6.040950E-6   -8.794298E-5   8.815022E-5   -1.760704E+2   -8.607043E+1   
4.822262E+3   1.100009E+2   1.100009E+2   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   -6.092721E-2   7.835579E-2   -8.870034E-5   -6.163141E-6   6.163141E-6   -8.870034E-5   8.891420E-5   -1.760253E+2   -8.602532E+1   
4.843962E+3   1.099716E+2   1.099716E+2   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   -6.320606E-2   8.043921E-2   -9.146615E-5   -5.839721E-6   5.839721E-6   -9.146615E-5   9.165238E-5   -1.763469E+2   -8.634687E+1   
4.865654E+3   1.100207E+2   1.100207E+2   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   -6.338861E-2   8.082516E-2   -9.183037E-5   -5.957023E-6   5.957023E-6   -9.183037E-5   9.202339E-5   -1.762884E+2   -8.628843E+1   
4.887374E+3   1.100416E+2   1.100416E+2   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   -6.362299E-2   8.291013E-2   -9.333320E-5   -7.146758E-6   7.146758E-6   -9.333320E-5   9.360642E-5   -1.756213E+2   -8.562126E+1   
4.909004E+3   1.100813E+2   1.100813E+2   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   -6.538583E-2   8.426891E-2   -9.530803E-5   -6.731244E-6   6.731244E-6   -9.530803E-5   9.554544E-5   -1.759601E+2   -8.596012E+1   
4.930681E+3   1.100441E+2   1.100441E+2   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   -6.727353E-2   8.618575E-2   -9.772351E-5   -6.588219E-6   6.588219E-6   -9.772351E-5   9.794533E-5   -1.761431E+2   -8.614313E+1   
4.952258E+3   1.100659E+2   1.100659E+2   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   -6.687930E-2   8.733008E-2   -9.822507E-5   -7.627930E-6   7.627930E-6   -9.822507E-5   9.852081E-5   -1.755595E+2   -8.555946E+1   
4.985312E+3   1.100086E+2   1.100086E+2   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   -6.584508E-2   8.672570E-2   -9.719204E-5   -7.997746E-6   7.997746E-6   -9.719204E-5   9.752055E-5   -1.752958E+2   -8.529584E+1   
5.007513E+3   1.100109E+2   1.100109E+2   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   -6.779632E-2   8.603205E-2   -9.794662E-5   -6.101061E-6   6.101061E-6   -9.794662E-5   9.813645E-5   -1.764357E+2   -8.643567E+1   
5.029810E+3   1.100124E+2   1.100124E+2   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   -6.742693E-2   8.686838E-2   -9.826293E-5   -6.921039E-6   6.921039E-6   -9.826293E-5   9.850637E-5   -1.759711E+2   -8.597109E+1   
5.052042E+3   1.100536E+2   1.100536E+2   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   -6.719099E-2   8.689290E-2   -9.813304E-5   -7.111580E-6   7.111580E-6   -9.813304E-5   9.839039E-5   -1.758551E+2   -8.585509E+1   
5.074311E+3   1.100388E+2   1.100388E+2   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   -6.629242E-2   8.766758E-2   -9.808204E-5   -8.282651E-6   8.282651E-6   -9.808204E-5   9.843114E-5   -1.751730E+2   -8.517304E+1   
5.096512E+3   1.100223E+2   1.100223E+2   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   -6.732323E-2   8.725186E-2   -9.844858E-5   -7.248447E-6   7.248447E-6   -9.844858E-5   9.871506E-5   -1.757891E+2   -8.578910E+1   
5.118774E+3   1.101074E+2   1.101074E+2   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   -6.613256E-2   8.715429E-2   -9.764891E-5   -8.065316E-6   8.065316E-6   -9.764891E-5   9.798142E-5   -1.752784E+2   -8.527837E+1   
5.141017E+3   1.099818E+2   1.099818E+2   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   -6.648937E-2   8.716718E-2   -9.787790E-5   -7.809840E-6   7.809840E-6   -9.787790E-5   9.818899E-5   -1.754379E+2   -8.543794E+1   
5.163303E+3   1.100301E+2   1.100301E+2   -3.100000E+1   -3.100000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   -6.690630E-2   8.719418E-2   -9.815325E-5   -7.519118E-6   7.519118E-6   -9.815325E-5   9.844083E-5   -1.756194E+2   -8.561936E+1   
5.184584E+3   1.100680E+2   1.100680E+2   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   -6.777789E-2   8.698433E-2   -9.855543E-5   -6.737271E-6   6.737271E-6   -9.855543E-5   9.878545E-5   -1.760893E+2   -8.608933E+1   
5.206864E+3   1.100353E+2   1.100353E+2   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   -6.784754E-2   8.690304E-2   -9.854555E-5   -6.632605E-6   6.632605E-6   -9.854555E-5   9.876850E-5   -1.761495E+2   -8.614952E+1   
5.229113E+3   1.100438E+2   1.100438E+2   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   -6.732015E-2   8.782125E-2   -9.881751E-5   -7.622976E-6   7.622976E-6   -9.881751E-5   9.911110E-5   -1.755888E+2   -8.558883E+1   
5.251354E+3   1.100183E+2   1.100183E+2   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   -6.657710E-2   8.767001E-2   -9.825962E-5   -8.073684E-6   8.073684E-6   -9.825962E-5   9.859076E-5   -1.753027E+2   -8.530274E+1   
5.273628E+3   1.100046E+2   1.100046E+2   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   -6.764628E-2   8.815384E-2   -9.923575E-5   -7.599200E-6   7.599200E-6   -9.923575E-5   9.952629E-5   -1.756210E+2   -8.562099E+1   
5.295873E+3   1.099921E+2   1.099921E+2   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.800000E+1   -1.800000E+1   -6.688359E-2   8.841678E-2   -9.893548E-5   -8.335208E-6   8.335208E-6   -9.893548E-5   9.928597E-5   -1.751843E+2   -8.518426E+1   
5.318113E+3   1.099983E+2   1.099983E+2   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   -6.792853E-2   8.776850E-2   -9.915929E-5   -7.138512E-6   7.138512E-6   -9.915929E-5   9.941591E-5   -1.758824E+2   -8.588236E+1   
5.340381E+3   1.099337E+2   1.099337E+2   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   -6.704189E-2   8.773353E-2   -9.858835E-5   -7.771442E-6   7.771442E-6   -9.858835E-5   9.889418E-5   -1.754929E+2   -8.549286E+1   
5.362658E+3   1.100403E+2   1.100403E+2   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   -6.762695E-2   8.823943E-2   -9.927955E-5   -7.669448E-6   7.669448E-6   -9.927955E-5   9.957534E-5   -1.755826E+2   -8.558261E+1   
5.384918E+3   1.100802E+2   1.100802E+2   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   -6.647096E-2   8.806271E-2   -9.844977E-5   -8.408925E-6   8.408925E-6   -9.844977E-5   9.880823E-5   -1.751180E+2   -8.511802E+1   
5.407159E+3   1.099943E+2   1.099943E+2   -1.000000E+1   -1.000000E+1   9.000000E+1   -8.000000E+0   -8.000000E+0   -6.713300E-2   8.855298E-2   -9.917837E-5   -8.239784E-6   8.239784E-6   -9.917837E-5   9.952007E-5   -1.752507E+2   -8.525075E+1   
5.429256E+3   1.100226E+2   1.100226E+2   -8.000000E+0   -8.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   -6.758124E-2   8.683431E-2   -9.833615E-5   -6.784630E-6   6.784630E-6   -9.833615E-5   9.856992E-5   -1.760532E+2   -8.605317E+1   
5.451327E+3   1.100338E+2   1.100338E+2   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   -6.801811E-2   8.871157E-2   -9.982889E-5   -7.688813E-6   7.688813E-6   -9.982889E-5   1.001245E-4   -1.755958E+2   -8.559578E+1   
5.473357E+3   1.100282E+2   1.100282E+2   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   -6.636818E-2   8.855142E-2   -9.870452E-5   -8.804451E-6   8.804451E-6   -9.870452E-5   9.909642E-5   -1.749027E+2   -8.490270E+1   
5.495400E+3   1.100221E+2   1.100221E+2   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   -6.823041E-2   8.793539E-2   -9.945462E-5   -7.024344E-6   7.024344E-6   -9.945462E-5   9.970237E-5   -1.759600E+2   -8.595999E+1   
5.517467E+3   1.099971E+2   1.099971E+2   0.000000E+0   0.000000E+0   9.000000E+1   0.000000E+0   0.000000E+0   -6.832706E-2   8.799001E-2   -9.954995E-5   -6.988571E-6   6.988571E-6   -9.954995E-5   9.979495E-5   -1.759843E+2   -8.598433E+1   
5.539445E+3   1.100053E+2   1.100053E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   -6.724348E-2   8.866557E-2   -9.932002E-5   -8.231679E-6   8.231679E-6   -9.932002E-5   9.966055E-5   -1.752621E+2   -8.526213E+1   
5.560920E+3   1.099797E+2   1.099797E+2   3.000000E+0   3.000000E+0   9.000000E+1   4.000000E+0   4.000000E+0   -6.675934E-2   8.785839E-2   -9.849499E-5   -8.062056E-6   8.062056E-6   -9.849499E-5   9.882438E-5   -1.753206E+2   -8.532063E+1   
5.582645E+3   1.100201E+2   1.100201E+2   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   -6.785581E-2   8.762921E-2   -9.902361E-5   -7.101237E-6   7.101237E-6   -9.902361E-5   9.927791E-5   -1.758982E+2   -8.589819E+1   
5.604165E+3   1.100744E+2   1.100744E+2   7.000000E+0   7.000000E+0   9.000000E+1   8.000000E+0   8.000000E+0   -6.755087E-2   8.737457E-2   -9.866924E-5   -7.160307E-6   7.160307E-6   -9.866924E-5   9.892871E-5   -1.758494E+2   -8.584939E+1   
5.625910E+3   1.100416E+2   1.100416E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   -6.764995E-2   8.807129E-2   -9.918426E-5   -7.542513E-6   7.542513E-6   -9.918426E-5   9.947064E-5   -1.756513E+2   -8.565129E+1   
5.647778E+3   1.099777E+2   1.099777E+2   1.000000E+1   1.000000E+1   9.000000E+1   1.100000E+1   1.100000E+1   -6.768341E-2   8.811272E-2   -9.923193E-5   -7.544860E-6   7.544860E-6   -9.923193E-5   9.951834E-5   -1.756520E+2   -8.565202E+1   
5.669713E+3   1.100610E+2   1.100610E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   -6.695201E-2   8.940462E-2   -9.962114E-5   -8.930428E-6   8.930428E-6   -9.962114E-5   1.000206E-4   -1.748775E+2   -8.487747E+1   
5.691548E+3   1.099982E+2   1.099982E+2   1.500000E+1   1.500000E+1   9.000000E+1   1.500000E+1   1.500000E+1   -6.768156E-2   8.820782E-2   -9.929273E-5   -7.608399E-6   7.608399E-6   -9.929273E-5   9.958380E-5   -1.756182E+2   -8.561822E+1   
5.713602E+3   1.100232E+2   1.100232E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   -6.706275E-2   8.914385E-2   -9.951977E-5   -8.678043E-6   8.678043E-6   -9.951977E-5   9.989742E-5   -1.750165E+2   -8.501646E+1   
5.735451E+3   1.100626E+2   1.100626E+2   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   -6.807795E-2   8.835233E-2   -9.963190E-5   -7.409691E-6   7.409691E-6   -9.963190E-5   9.990706E-5   -1.757467E+2   -8.574671E+1   
5.757420E+3   1.100296E+2   1.100296E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   -6.805340E-2   8.759731E-2   -9.912500E-5   -6.934237E-6   6.934237E-6   -9.912500E-5   9.936724E-5   -1.759984E+2   -8.599842E+1   
5.779343E+3   1.100723E+2   1.100723E+2   2.200000E+1   2.200000E+1   9.000000E+1   2.300000E+1   2.300000E+1   -6.749842E-2   8.845417E-2   -9.933994E-5   -7.904916E-6   7.904916E-6   -9.933994E-5   9.965396E-5   -1.754503E+2   -8.545031E+1   
5.801234E+3   1.100461E+2   1.100461E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   -6.736434E-2   8.866618E-2   -9.939513E-5   -8.142686E-6   8.142686E-6   -9.939513E-5   9.972811E-5   -1.753167E+2   -8.531665E+1   
5.823113E+3   1.100486E+2   1.100486E+2   2.600000E+1   2.600000E+1   9.000000E+1   2.700000E+1   2.700000E+1   -6.830406E-2   8.909845E-2   -1.002576E-4   -7.730249E-6   7.730249E-6   -1.002576E-4   1.005552E-4   -1.755910E+2   -8.559100E+1   
5.845003E+3   1.100038E+2   1.100038E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   -6.804757E-2   8.801149E-2   -9.939114E-5   -7.209328E-6   7.209328E-6   -9.939114E-5   9.965226E-5   -1.758513E+2   -8.585132E+1   
5.866880E+3   1.100386E+2   1.100386E+2   3.100000E+1   3.100000E+1   9.000000E+1   3.100000E+1   3.100000E+1   -6.787945E-2   8.889932E-2   -9.986544E-5   -7.914114E-6   7.914114E-6   -9.986544E-5   1.001785E-4   -1.754689E+2   -8.546891E+1   
5.888918E+3   1.100385E+2   1.100385E+2   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   -6.814481E-2   8.801269E-2   -9.945205E-5   -7.138194E-6   7.138194E-6   -9.945205E-5   9.970789E-5   -1.758946E+2   -8.589462E+1   
5.910847E+3   1.100471E+2   1.100471E+2   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   -6.851543E-2   8.941997E-2   -1.005977E-4   -7.784109E-6   7.784109E-6   -1.005977E-4   1.008984E-4   -1.755754E+2   -8.557535E+1   
5.932822E+3   1.099929E+2   1.099929E+2   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   -6.758124E-2   8.913926E-2   -9.983734E-5   -8.291546E-6   8.291546E-6   -9.983734E-5   1.001811E-4   -1.752524E+2   -8.525245E+1   
5.954781E+3   1.100115E+2   1.100115E+2   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   -6.722597E-2   8.929018E-2   -9.971598E-5   -8.652981E-6   8.652981E-6   -9.971598E-5   1.000907E-4   -1.750405E+2   -8.504051E+1   
5.976655E+3   1.099770E+2   1.099770E+2   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   -6.801687E-2   8.983105E-2   -1.005572E-4   -8.421609E-6   8.421609E-6   -1.005572E-4   1.009093E-4   -1.752127E+2   -8.521268E+1   
5.998520E+3   1.099748E+2   1.099748E+2   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   -6.778526E-2   9.004183E-2   -1.005513E-4   -8.730722E-6   8.730722E-6   -1.005513E-4   1.009296E-4   -1.750375E+2   -8.503754E+1   
6.020400E+3   1.100135E+2   1.100135E+2   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   -6.734809E-2   9.013542E-2   -1.003420E-4   -9.115249E-6   9.115249E-6   -1.003420E-4   1.007552E-4   -1.748094E+2   -8.480939E+1   
6.042341E+3   1.100658E+2   1.100658E+2   4.600000E+1   4.600000E+1   9.000000E+1   4.700000E+1   4.700000E+1   -6.860224E-2   8.915950E-2   -1.004818E-4   -7.549616E-6   7.549616E-6   -1.004818E-4   1.007650E-4   -1.757032E+2   -8.570320E+1   
6.064210E+3   1.100538E+2   1.100538E+2   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   -6.802578E-2   8.938529E-2   -1.002724E-4   -8.123601E-6   8.123601E-6   -1.002724E-4   1.006009E-4   -1.753683E+2   -8.536828E+1   
6.098072E+3   1.099862E+2   1.099862E+2   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   -6.909833E-2   9.034771E-2   -1.015623E-4   -7.959515E-6   7.959515E-6   -1.015623E-4   1.018737E-4   -1.755188E+2   -8.551885E+1   
6.120411E+3   1.100018E+2   1.100018E+2   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   -7.069059E-2   9.188111E-2   -1.035454E-4   -7.784319E-6   7.784319E-6   -1.035454E-4   1.038376E-4   -1.757007E+2   -8.570072E+1   
6.142794E+3   1.099885E+2   1.099885E+2   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   -7.093633E-2   9.353326E-2   -1.047734E-4   -8.682688E-6   8.682688E-6   -1.047734E-4   1.051325E-4   -1.752627E+2   -8.526266E+1   
6.165123E+3   1.100451E+2   1.100451E+2   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   -7.306025E-2   9.434632E-2   -1.066160E-4   -7.643330E-6   7.643330E-6   -1.066160E-4   1.068896E-4   -1.758995E+2   -8.589947E+1   
6.187743E+3   1.100131E+2   1.100131E+2   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   -7.451355E-2   9.491790E-2   -1.078868E-4   -6.942110E-6   6.942110E-6   -1.078868E-4   1.081099E-4   -1.763183E+2   -8.631831E+1   
6.210032E+3   1.100302E+2   1.100302E+2   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   -7.445922E-2   9.758558E-2   -1.095906E-4   -8.726349E-6   8.726349E-6   -1.095906E-4   1.099375E-4   -1.754473E+2   -8.544733E+1   
6.232220E+3   1.099610E+2   1.099610E+2   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   -7.492586E-2   9.965092E-2   -1.112243E-4   -9.731465E-6   9.731465E-6   -1.112243E-4   1.116492E-4   -1.749997E+2   -8.499969E+1   
6.255102E+3   1.100622E+2   1.100622E+2   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   -7.630795E-2   1.002400E-1   -1.124624E-4   -9.094322E-6   9.094322E-6   -1.124624E-4   1.128295E-4   -1.753768E+2   -8.537681E+1   
6.277286E+3   1.099748E+2   1.099748E+2   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   -7.636746E-2   1.021706E-1   -1.137566E-4   -1.031251E-5   1.031251E-5   -1.137566E-4   1.142231E-4   -1.748201E+2   -8.482006E+1   
6.299927E+3   1.100038E+2   1.100038E+2   5.480000E+2   5.480000E+2   9.000000E+1   5.480000E+2   5.480000E+2   -7.827110E-2   1.030496E-1   -1.155059E-4   -9.479157E-6   9.479157E-6   -1.155059E-4   1.158943E-4   -1.753085E+2   -8.530846E+1   
6.323258E+3   1.100150E+2   1.100150E+2   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   -7.901753E-2   1.041792E-1   -1.167031E-4   -9.665584E-6   9.665584E-6   -1.167031E-4   1.171027E-4   -1.752655E+2   -8.526546E+1   
6.345887E+3   1.100559E+2   1.100559E+2   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   -8.020576E-2   1.053766E-1   -1.182176E-4   -9.569559E-6   9.569559E-6   -1.182176E-4   1.186043E-4   -1.753721E+2   -8.537207E+1   
6.368469E+3   1.100170E+2   1.100170E+2   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   -8.077608E-2   1.079598E-1   -1.202526E-4   -1.083657E-5   1.083657E-5   -1.202526E-4   1.207399E-4   -1.748507E+2   -8.485070E+1   
6.391854E+3   1.099909E+2   1.099909E+2   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   -8.046068E-2   1.090986E-1   -1.207993E-4   -1.181438E-5   1.181438E-5   -1.207993E-4   1.213757E-4   -1.744141E+2   -8.441414E+1   
6.414479E+3   1.100475E+2   1.100475E+2   7.970000E+2   7.970000E+2   9.000000E+1   7.980000E+2   7.980000E+2   -8.224745E-2   1.109096E-1   -1.230835E-4   -1.167679E-5   1.167679E-5   -1.230835E-4   1.236361E-4   -1.745806E+2   -8.458063E+1   
6.437047E+3   1.100369E+2   1.100369E+2   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   -8.297609E-2   1.108375E-1   -1.234870E-4   -1.109074E-5   1.109074E-5   -1.234870E-4   1.239840E-4   -1.748679E+2   -8.486786E+1   
6.460389E+3   1.101348E+2   1.101348E+2   8.970000E+2   8.970000E+2   9.000000E+1   8.980000E+2   8.980000E+2   -8.297455E-2   1.135241E-1   -1.252358E-4   -1.284828E-5   1.284828E-5   -1.252358E-4   1.258931E-4   -1.741424E+2   -8.414236E+1   
6.483032E+3   1.099898E+2   1.099898E+2   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   -8.409557E-2   1.149826E-1   -1.268788E-4   -1.297267E-5   1.297267E-5   -1.268788E-4   1.275402E-4   -1.741621E+2   -8.416210E+1   
6.505602E+3   1.100505E+2   1.100505E+2   9.980000E+2   9.980000E+2   9.000000E+1   9.980000E+2   9.980000E+2   -8.562126E-2   1.163733E-1   -1.287277E-4   -1.275341E-5   1.275341E-5   -1.287277E-4   1.293580E-4   -1.743420E+2   -8.434201E+1   
6.529194E+3   1.100375E+2   1.100375E+2   1.048000E+3   1.048000E+3   9.000000E+1   1.048000E+3   1.048000E+3   -8.692849E-2   1.172268E-1   -1.300918E-4   -1.234454E-5   1.234454E-5   -1.300918E-4   1.306762E-4   -1.745794E+2   -8.457938E+1   
6.552016E+3   1.099988E+2   1.099988E+2   1.097000E+3   1.097000E+3   9.000000E+1   1.098000E+3   1.098000E+3   -8.789765E-2   1.181591E-1   -1.312982E-4   -1.223726E-5   1.223726E-5   -1.312982E-4   1.318672E-4   -1.746753E+2   -8.467530E+1   
6.574848E+3   1.100121E+2   1.100121E+2   1.148000E+3   1.148000E+3   9.000000E+1   1.148000E+3   1.148000E+3   -8.828206E-2   1.207144E-1   -1.332001E-4   -1.362350E-5   1.362350E-5   -1.332001E-4   1.338950E-4   -1.741602E+2   -8.416018E+1   
6.598390E+3   1.100318E+2   1.100318E+2   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   -8.820169E-2   1.213154E-1   -1.335418E-4   -1.407587E-5   1.407587E-5   -1.335418E-4   1.342816E-4   -1.739830E+2   -8.398300E+1   
6.621231E+3   1.100368E+2   1.100368E+2   1.248000E+3   1.248000E+3   9.000000E+1   1.248000E+3   1.248000E+3   -8.790687E-2   1.237869E-1   -1.349692E-4   -1.590974E-5   1.590974E-5   -1.349692E-4   1.359037E-4   -1.732772E+2   -8.327718E+1   
6.644066E+3   1.100151E+2   1.100151E+2   1.298000E+3   1.298000E+3   9.000000E+1   1.298000E+3   1.298000E+3   -9.019127E-2   1.246438E-1   -1.369396E-4   -1.478033E-5   1.478033E-5   -1.369396E-4   1.377350E-4   -1.738397E+2   -8.383973E+1   
6.667340E+3   1.100313E+2   1.100313E+2   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   -9.084687E-2   1.259645E-1   -1.382051E-4   -1.515888E-5   1.515888E-5   -1.382051E-4   1.390340E-4   -1.737406E+2   -8.374060E+1   
6.689931E+3   1.100579E+2   1.100579E+2   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   -9.163383E-2   1.277267E-1   -1.398394E-4   -1.572891E-5   1.572891E-5   -1.398394E-4   1.407212E-4   -1.735824E+2   -8.358244E+1   
6.712964E+3   1.100755E+2   1.100755E+2   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   -9.432303E-2   1.283928E-1   -1.419358E-4   -1.417533E-5   1.417533E-5   -1.419358E-4   1.426419E-4   -1.742967E+2   -8.429670E+1   
6.736052E+3   1.099900E+2   1.099900E+2   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   -9.466664E-2   1.314592E-1   -1.441453E-4   -1.592592E-5   1.592592E-5   -1.441453E-4   1.450224E-4   -1.736952E+2   -8.369524E+1   
6.758677E+3   1.099660E+2   1.099660E+2   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   -9.603501E-2   1.316061E-1   -1.450870E-4   -1.500990E-5   1.500990E-5   -1.450870E-4   1.458614E-4   -1.740935E+2   -8.409351E+1   
6.781211E+3   1.100811E+2   1.100811E+2   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   -9.682867E-2   1.336715E-1   -1.469228E-4   -1.577314E-5   1.577314E-5   -1.469228E-4   1.477671E-4   -1.738724E+2   -8.387239E+1   
6.804245E+3   1.100106E+2   1.100106E+2   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   -9.536735E-2   1.348624E-1   -1.467950E-4   -1.763260E-5   1.763260E-5   -1.467950E-4   1.478502E-4   -1.731506E+2   -8.315061E+1   
6.826765E+3   1.100658E+2   1.100658E+2   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   -9.767516E-2   1.363486E-1   -1.491897E-4   -1.689725E-5   1.689725E-5   -1.491897E-4   1.501436E-4   -1.735382E+2   -8.353821E+1   
6.849301E+3   1.099833E+2   1.099833E+2   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   -9.962977E-2   1.379960E-1   -1.514711E-4   -1.652862E-5   1.652862E-5   -1.514711E-4   1.523703E-4   -1.737725E+2   -8.377249E+1   
6.872122E+3   1.100156E+2   1.100156E+2   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   -9.677285E-2   1.396340E-1   -1.507716E-4   -1.971255E-5   1.971255E-5   -1.507716E-4   1.520548E-4   -1.725511E+2   -8.255115E+1   
6.894667E+3   1.099773E+2   1.099773E+2   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   -1.007005E-1   1.403586E-1   -1.536718E-4   -1.728131E-5   1.728131E-5   -1.536718E-4   1.546405E-4   -1.735837E+2   -8.358371E+1   
6.917211E+3   1.100680E+2   1.100680E+2   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   -1.009962E-1   1.412907E-1   -1.544617E-4   -1.767189E-5   1.767189E-5   -1.544617E-4   1.554693E-4   -1.734732E+2   -8.347319E+1   
6.940004E+3   1.100051E+2   1.100051E+2   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   -1.013316E-1   1.432725E-1   -1.559598E-4   -1.871956E-5   1.871956E-5   -1.559598E-4   1.570792E-4   -1.731556E+2   -8.315564E+1   
6.962541E+3   1.100615E+2   1.100615E+2   1.999000E+3   1.999000E+3   9.000000E+1   1.999000E+3   1.999000E+3   -1.030965E-1   1.463445E-1   -1.590517E-4   -1.942249E-5   1.942249E-5   -1.590517E-4   1.602332E-4   -1.730378E+2   -8.303784E+1   
7.000448E+3   1.099853E+2   1.099853E+2   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   -1.118548E-1   1.600510E-1   -1.733934E-4   -2.190554E-5   2.190554E-5   -1.733934E-4   1.747717E-4   -1.727997E+2   -8.279972E+1   
7.027284E+3   1.099497E+2   1.099497E+2   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   -1.229770E-1   1.774274E-1   -1.915867E-4   -2.503946E-5   2.503946E-5   -1.915867E-4   1.932161E-4   -1.725539E+2   -8.255392E+1   
7.052924E+3   1.100076E+2   1.100076E+2   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -1.314273E-1   1.923649E-1   -2.065397E-4   -2.855505E-5   2.855505E-5   -2.065397E-4   2.085043E-4   -1.721285E+2   -8.212850E+1   
7.078859E+3   1.099584E+2   1.099584E+2   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -1.412075E-1   2.061096E-1   -2.215381E-4   -3.030716E-5   3.030716E-5   -2.215381E-4   2.236015E-4   -1.722101E+2   -8.221010E+1   
7.105558E+3   1.100017E+2   1.100017E+2   4.498000E+3   4.498000E+3   9.000000E+1   4.499000E+3   4.499000E+3   -1.445626E-1   2.152360E-1   -2.295563E-4   -3.379226E-5   3.379226E-5   -2.295563E-4   2.320302E-4   -1.716258E+2   -8.162581E+1   
7.131764E+3   1.100076E+2   1.100076E+2   4.998000E+3   4.998000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -1.375346E-1   2.106204E-1   -2.222051E-4   -3.597279E-5   3.597279E-5   -2.222051E-4   2.250981E-4   -1.708042E+2   -8.080417E+1   
7.157410E+3   1.099784E+2   1.099784E+2   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -1.258933E-1   1.990564E-1   -2.074765E-4   -3.702285E-5   3.702285E-5   -2.074765E-4   2.107539E-4   -1.698824E+2   -7.988243E+1   
7.183863E+3   1.100375E+2   1.100375E+2   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -1.070520E-1   1.793200E-1   -1.829738E-4   -3.805540E-5   3.805540E-5   -1.829738E-4   1.868893E-4   -1.682510E+2   -7.825096E+1   
7.209808E+3   1.099850E+2   1.099850E+2   6.498000E+3   6.498000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -8.959240E-2   1.628711E-1   -1.614664E-4   -4.021518E-5   4.021518E-5   -1.614664E-4   1.663991E-4   -1.660143E+2   -7.601434E+1   
7.235973E+3   1.099489E+2   1.099489E+2   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -8.259475E-2   1.538060E-1   -1.512361E-4   -3.946434E-5   3.946434E-5   -1.512361E-4   1.563003E-4   -1.653751E+2   -7.537507E+1   
7.261622E+3   1.100128E+2   1.100128E+2   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -7.941883E-2   1.520747E-1   -1.481451E-4   -4.068153E-5   4.068153E-5   -1.481451E-4   1.536293E-4   -1.646447E+2   -7.464474E+1   
7.287521E+3   1.100283E+2   1.100283E+2   7.998000E+3   7.998000E+3   9.000000E+1   8.000000E+3   8.000000E+3   -8.132861E-2   1.597053E-1   -1.542955E-4   -4.425762E-5   4.425762E-5   -1.542955E-4   1.605174E-4   -1.639952E+2   -7.399516E+1   
7.313962E+3   1.100159E+2   1.100159E+2   8.497000E+3   8.497000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -8.956084E-2   1.745488E-1   -1.690525E-4   -4.787309E-5   4.787309E-5   -1.690525E-4   1.757002E-4   -1.641887E+2   -7.418868E+1   
7.340614E+3   1.100563E+2   1.100563E+2   8.998000E+3   8.998000E+3   9.000000E+1   8.999000E+3   8.999000E+3   -9.458501E-2   1.842985E-1   -1.785086E-4   -5.053118E-5   5.053118E-5   -1.785086E-4   1.855228E-4   -1.641945E+2   -7.419455E+1   
7.366971E+3   1.100536E+2   1.100536E+2   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -1.056589E-1   2.033880E-1   -1.977877E-4   -5.482078E-5   5.482078E-5   -1.977877E-4   2.052445E-4   -1.645082E+2   -7.450823E+1   
7.392902E+3   1.100012E+2   1.100012E+2   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -1.211479E-1   2.215005E-1   -2.191602E-4   -5.520600E-5   5.520600E-5   -2.191602E-4   2.260064E-4   -1.658615E+2   -7.586146E+1   
@@END Data.
@Time at end of measurement: 12:55:33
@NO Instrument  Changes.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -9499.000      -9998.000      249.500        Coercive Field: Field at which M//H changes sign
Ms  emu                                 2.738E-4       -3.261E-4      3.000E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -9.955E-5      1.303E-4       1.149E-4       Remanent Magnetization: M at H=0        
S                                       0.364          0.400          0.382          Squareness: Mr/Ms                       
S*                                      1.331          1.342          1.336          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
