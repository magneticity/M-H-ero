@Filename: c:\vsm-lv\Will\data\AJA335e-FePtFeRh_1030nm_Tann_6\AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_RT.VHD
@Measurement Controlfilename: c:\vsm-lv\Will\Recipes\10kOe OoP loop.VHC
@Signal Manipulation filename: c:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA335e-FePtFeRh_1030nm_Tann_600C
@Date: 05 November 2019    (2019-05-11)
@Time: 10:43:37
@Test ID: AJA335e_FePt_FeRh_Pt_600deg_annealed_OoP_RT
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 90.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Applied Field to 10000.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Auto Range Signal to 12.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 5
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 5.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 10000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To: 50.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: 50.0000 [Oe] To: -50.0000 [Oe] Min Stepsize/Sweeprate =  2.0000 [Oe] Max Stepsize/Sweeprate =  2.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -50.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -10000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 4 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 20 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.706
@Y Coils Correction Factor: 0.964
@Sample Shape Correction Factor: 0.919
@Coil Angle Alpha: 42.300
@Coil Angle Beta: -47.320
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
15000.000000   1.000000
15249.000000   1.000524
15499.000000   1.000702
15750.000000   1.001233
16000.000000   1.001406
16250.000000   1.001585
16499.000000   1.001758
16749.000000   1.001937
16999.000000   1.002110
17249.000000   1.001937
17499.000000   1.002289
17749.000000   1.002289
17999.000000   1.002289
18249.000000   1.002462
18499.000000   1.002462
18748.000000   1.002462
18999.000000   1.002462
19249.000000   1.002462
19499.000000   1.002642
19749.000000   1.002642
19999.000000   1.002462
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = No
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 25 October 2019  12:02:56
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 5
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 10:43:37
@@Data
New Section: Section 0: 
2.964500E+1   2.082980E+1   2.082980E+1   9.999000E+3   9.999000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -2.069821E-1   2.830499E-1   -3.123134E-4   -3.195962E-5   3.195962E-5   -3.123134E-4   3.139444E-4   -1.741572E+2   -8.415715E+1   
5.498300E+1   2.082760E+1   2.082760E+1   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -1.852632E-1   2.587689E-1   -2.830718E-4   -3.214942E-5   3.214942E-5   -2.830718E-4   2.848916E-4   -1.735205E+2   -8.352049E+1   
8.010100E+1   2.079849E+1   2.079849E+1   8.998000E+3   8.998000E+3   9.000000E+1   8.998000E+3   8.998000E+3   -1.619025E-1   2.331472E-1   -2.519420E-4   -3.267693E-5   3.267693E-5   -2.519420E-4   2.540523E-4   -1.726100E+2   -8.260998E+1   
1.051800E+2   2.079910E+1   2.079910E+1   8.498000E+3   8.498000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -1.405577E-1   2.056555E-1   -2.208406E-4   -3.049091E-5   3.049091E-5   -2.208406E-4   2.229356E-4   -1.721390E+2   -8.213901E+1   
1.309180E+2   2.079370E+1   2.079370E+1   7.999000E+3   7.999000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -1.227033E-1   1.834416E-1   -1.953345E-4   -2.917374E-5   2.917374E-5   -1.953345E-4   1.975011E-4   -1.715055E+2   -8.150551E+1   
1.563230E+2   2.078640E+1   2.078640E+1   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -1.060770E-1   1.616776E-1   -1.708807E-4   -2.724240E-5   2.724240E-5   -1.708807E-4   1.730386E-4   -1.709419E+2   -8.094193E+1   
1.816430E+2   2.079049E+1   2.079049E+1   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -8.921199E-2   1.403326E-1   -1.465521E-4   -2.576150E-5   2.576150E-5   -1.465521E-4   1.487991E-4   -1.700302E+2   -8.003018E+1   
2.072290E+2   2.076660E+1   2.076660E+1   6.498000E+3   6.498000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -7.202790E-2   1.173633E-1   -1.209685E-4   -2.345474E-5   2.345474E-5   -1.209685E-4   1.232213E-4   -1.690270E+2   -7.902700E+1   
2.323130E+2   2.076071E+1   2.076071E+1   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -5.835167E-2   9.942569E-2   -1.008306E-4   -2.184300E-5   2.184300E-5   -1.008306E-4   1.031694E-4   -1.677769E+2   -7.777685E+1   
2.576950E+2   2.075302E+1   2.075302E+1   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -3.981265E-2   7.653804E-2   -7.446245E-5   -2.059173E-5   2.059173E-5   -7.446245E-5   7.725721E-5   -1.645418E+2   -7.454183E+1   
2.830830E+2   2.072790E+1   2.072790E+1   4.998000E+3   4.998000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -2.562377E-2   5.633760E-2   -5.253390E-5   -1.787979E-5   1.787979E-5   -5.253390E-5   5.549322E-5   -1.612041E+2   -7.120411E+1   
3.082590E+2   2.071060E+1   2.071060E+1   4.498000E+3   4.498000E+3   9.000000E+1   4.498000E+3   4.498000E+3   -1.178857E-2   3.840387E-2   -3.230028E-5   -1.638817E-5   1.638817E-5   -3.230028E-5   3.621989E-5   -1.530982E+2   -6.309816E+1   
3.341070E+2   2.070541E+1   2.070541E+1   3.999000E+3   3.999000E+3   9.000000E+1   3.999000E+3   3.999000E+3   9.961616E-4   2.065736E-2   -1.283805E-5   -1.424199E-5   1.424199E-5   -1.283805E-5   1.917420E-5   -1.320322E+2   -4.203220E+1   
3.595130E+2   2.070910E+1   2.070910E+1   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   1.627697E-2   -5.556044E-4   1.042504E-5   -1.167571E-5   1.167571E-5   1.042504E-5   1.565260E-5   -4.823889E+1   4.176111E+1   
3.843890E+2   2.069171E+1   2.069171E+1   2.998000E+3   2.998000E+3   9.000000E+1   2.998000E+3   2.998000E+3   2.864601E-2   -1.804563E-2   2.946323E-5   -9.389753E-6   9.389753E-6   2.946323E-5   3.092328E-5   -1.767676E+1   7.232324E+1   
4.098010E+2   2.067410E+1   2.067410E+1   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   4.355033E-2   -3.750739E-2   5.135302E-5   -7.689902E-6   7.689902E-6   5.135302E-5   5.192559E-5   -8.516525E+0   8.148348E+1   
4.356020E+2   2.067831E+1   2.067831E+1   1.999000E+3   1.999000E+3   9.000000E+1   1.999000E+3   1.999000E+3   5.758992E-2   -5.796912E-2   7.335945E-5   -4.696720E-6   4.696720E-6   7.335945E-5   7.350965E-5   -3.663270E+0   8.633673E+1   
4.694650E+2   2.067150E+1   2.067150E+1   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   5.950276E-2   -5.840968E-2   7.482899E-5   -5.823490E-6   5.823490E-6   7.482899E-5   7.505526E-5   -4.450016E+0   8.554998E+1   
4.917750E+2   2.066241E+1   2.066241E+1   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   6.115088E-2   -6.241485E-2   7.845646E-5   -4.424023E-6   4.424023E-6   7.845646E-5   7.858110E-5   -3.227391E+0   8.677261E+1   
5.140450E+2   2.064691E+1   2.064691E+1   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   6.253724E-2   -6.325331E-2   7.985966E-5   -4.901260E-6   4.901260E-6   7.985966E-5   8.000992E-5   -3.512032E+0   8.648797E+1   
5.362970E+2   2.063009E+1   2.063009E+1   1.799000E+3   1.799000E+3   9.000000E+1   1.799000E+3   1.799000E+3   6.407367E-2   -6.603747E-2   8.262284E-5   -4.217442E-6   4.217442E-6   8.262284E-5   8.273041E-5   -2.922098E+0   8.707790E+1   
5.585450E+2   2.061880E+1   2.061880E+1   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   6.441236E-2   -6.655748E-2   8.317091E-5   -4.127989E-6   4.127989E-6   8.317091E-5   8.327329E-5   -2.841407E+0   8.715859E+1   
5.808230E+2   2.061920E+1   2.061920E+1   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   6.773187E-2   -6.870135E-2   8.661947E-5   -5.181597E-6   5.181597E-6   8.661947E-5   8.677432E-5   -3.423367E+0   8.657663E+1   
6.031390E+2   2.062081E+1   2.062081E+1   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   6.891333E-2   -7.183953E-2   8.939377E-5   -4.003783E-6   4.003783E-6   8.939377E-5   8.948338E-5   -2.564459E+0   8.743554E+1   
6.253580E+2   2.061929E+1   2.061929E+1   1.599000E+3   1.599000E+3   9.000000E+1   1.599000E+3   1.599000E+3   6.905997E-2   -7.269546E-2   9.004189E-5   -3.552665E-6   3.552665E-6   9.004189E-5   9.011195E-5   -2.259473E+0   8.774053E+1   
6.476460E+2   2.060500E+1   2.060500E+1   1.549000E+3   1.549000E+3   9.000000E+1   1.549000E+3   1.549000E+3   7.144591E-2   -7.498813E-2   9.301018E-5   -3.818491E-6   3.818491E-6   9.301018E-5   9.308853E-5   -2.350932E+0   8.764907E+1   
6.698870E+2   2.059011E+1   2.059011E+1   1.499000E+3   1.499000E+3   9.000000E+1   1.499000E+3   1.499000E+3   7.259822E-2   -7.728847E-2   9.522078E-5   -3.166877E-6   3.166877E-6   9.522078E-5   9.527343E-5   -1.904856E+0   8.809514E+1   
6.921680E+2   2.059100E+1   2.059100E+1   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   7.371063E-2   -7.862698E-2   9.678028E-5   -3.114574E-6   3.114574E-6   9.678028E-5   9.683039E-5   -1.843251E+0   8.815675E+1   
7.144420E+2   2.058611E+1   2.058611E+1   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   7.552134E-2   -8.015054E-2   9.889202E-5   -3.457769E-6   3.457769E-6   9.889202E-5   9.895245E-5   -2.002537E+0   8.799746E+1   
7.364810E+2   2.057571E+1   2.057571E+1   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   7.668284E-2   -8.358260E-2   1.018454E-4   -2.073068E-6   2.073068E-6   1.018454E-4   1.018665E-4   -1.166098E+0   8.883390E+1   
7.586780E+2   2.058709E+1   2.058709E+1   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   7.808612E-2   -8.433395E-2   1.032023E-4   -2.619762E-6   2.619762E-6   1.032023E-4   1.032355E-4   -1.454125E+0   8.854587E+1   
7.809480E+2   2.056179E+1   2.056179E+1   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   7.960628E-2   -8.538227E-2   1.048249E-4   -3.058759E-6   3.058759E-6   1.048249E-4   1.048695E-4   -1.671399E+0   8.832860E+1   
8.032210E+2   2.056680E+1   2.056680E+1   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   8.091076E-2   -8.844465E-2   1.076259E-4   -2.021494E-6   2.021494E-6   1.076259E-4   1.076449E-4   -1.076037E+0   8.892396E+1   
8.255370E+2   2.055139E+1   2.055139E+1   1.148000E+3   1.148000E+3   9.000000E+1   1.149000E+3   1.149000E+3   8.189465E-2   -9.006456E-2   1.092892E-4   -1.690163E-6   1.690163E-6   1.092892E-4   1.093023E-4   -8.860114E-1   8.911399E+1   
8.477670E+2   2.055111E+1   2.055111E+1   1.098000E+3   1.098000E+3   9.000000E+1   1.099000E+3   1.099000E+3   8.322458E-2   -9.143010E-2   1.110008E-4   -1.781069E-6   1.781069E-6   1.110008E-4   1.110151E-4   -9.192638E-1   8.908074E+1   
8.700510E+2   2.052761E+1   2.052761E+1   1.048000E+3   1.048000E+3   9.000000E+1   1.048000E+3   1.048000E+3   8.563844E-2   -9.375630E-2   1.140082E-4   -2.045627E-6   2.045627E-6   1.140082E-4   1.140265E-4   -1.027937E+0   8.897206E+1   
8.922330E+2   2.052029E+1   2.052029E+1   9.980000E+2   9.980000E+2   9.000000E+1   9.990000E+2   9.990000E+2   8.689750E-2   -9.624977E-2   1.164106E-4   -1.346706E-6   1.346706E-6   1.164106E-4   1.164183E-4   -6.628020E-1   8.933720E+1   
9.140650E+2   2.050729E+1   2.050729E+1   9.480000E+2   9.480000E+2   9.000000E+1   9.480000E+2   9.480000E+2   8.724817E-2   -9.748496E-2   1.174318E-4   -7.985441E-7   7.985441E-7   1.174318E-4   1.174345E-4   -3.896091E-1   8.961039E+1   
9.358840E+2   2.050881E+1   2.050881E+1   8.980000E+2   8.980000E+2   9.000000E+1   8.980000E+2   8.980000E+2   8.801546E-2   -9.891584E-2   1.188381E-4   -4.305874E-7   4.305874E-7   1.188381E-4   1.188389E-4   -2.075995E-1   8.979240E+1   
9.577600E+2   2.050302E+1   2.050302E+1   8.480000E+2   8.480000E+2   9.000000E+1   8.480000E+2   8.480000E+2   8.878183E-2   -1.007541E-1   1.205092E-4   2.044148E-7   -2.044148E-7   1.205092E-4   1.205094E-4   9.718838E-2   9.009719E+1   
9.796460E+2   2.048019E+1   2.048019E+1   7.980000E+2   7.980000E+2   9.000000E+1   7.990000E+2   7.990000E+2   9.130184E-2   -1.017951E-1   1.227451E-4   -9.789121E-7   9.789121E-7   1.227451E-4   1.227490E-4   -4.569333E-1   8.954307E+1   
1.001525E+3   2.048330E+1   2.048330E+1   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   9.153075E-2   -1.046243E-1   1.247293E-4   7.014548E-7   -7.014548E-7   1.247293E-4   1.247313E-4   3.222176E-1   9.032222E+1   
1.023394E+3   2.046801E+1   2.046801E+1   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   9.277577E-2   -1.054981E-1   1.260681E-4   3.518356E-7   -3.518356E-7   1.260681E-4   1.260686E-4   1.599028E-1   9.015990E+1   
1.045212E+3   2.045419E+1   2.045419E+1   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   9.407294E-2   -1.066654E-1   1.276304E-4   1.555761E-7   -1.555761E-7   1.276304E-4   1.276305E-4   6.984113E-2   9.006984E+1   
1.067092E+3   2.046740E+1   2.046740E+1   5.980000E+2   5.980000E+2   9.000000E+1   5.990000E+2   5.990000E+2   9.694556E-2   -1.080116E-1   1.302831E-4   -1.088988E-6   1.088988E-6   1.302831E-4   1.302877E-4   -4.789029E-1   8.952110E+1   
1.088983E+3   2.045641E+1   2.045641E+1   5.480000E+2   5.480000E+2   9.000000E+1   5.480000E+2   5.480000E+2   9.636293E-2   -1.106786E-1   1.316599E-4   1.085516E-6   -1.085516E-6   1.316599E-4   1.316643E-4   4.723844E-1   9.047238E+1   
1.110853E+3   2.044781E+1   2.044781E+1   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   9.701705E-2   -1.132603E-1   1.337457E-4   2.289532E-6   -2.289532E-6   1.337457E-4   1.337653E-4   9.807249E-1   9.098072E+1   
1.132697E+3   2.044000E+1   2.044000E+1   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   9.864279E-2   -1.148939E-1   1.358148E-4   2.155127E-6   -2.155127E-6   1.358148E-4   1.358319E-4   9.091007E-1   9.090910E+1   
1.154587E+3   2.043270E+1   2.043270E+1   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   9.950703E-2   -1.158517E-1   1.369729E-4   2.142091E-6   -2.142091E-6   1.369729E-4   1.369896E-4   8.959640E-1   9.089596E+1   
1.176459E+3   2.043740E+1   2.043740E+1   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   1.009649E-1   -1.179204E-1   1.392216E-4   2.416257E-6   -2.416257E-6   1.392216E-4   1.392425E-4   9.942959E-1   9.099430E+1   
1.198293E+3   2.042370E+1   2.042370E+1   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   1.032453E-1   -1.191209E-1   1.414133E-4   1.514432E-6   -1.514432E-6   1.414133E-4   1.414214E-4   6.135723E-1   9.061357E+1   
1.220219E+3   2.043170E+1   2.043170E+1   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   1.029437E-1   -1.209531E-1   1.424201E-4   2.935322E-6   -2.935322E-6   1.424201E-4   1.424503E-4   1.180716E+0   9.118072E+1   
1.242046E+3   2.042629E+1   2.042629E+1   1.990000E+2   1.990000E+2   9.000000E+1   1.990000E+2   1.990000E+2   1.043826E-1   -1.213654E-1   1.435782E-4   2.140660E-6   -2.140660E-6   1.435782E-4   1.435942E-4   8.541806E-1   9.085418E+1   
1.263930E+3   2.042111E+1   2.042111E+1   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   1.054263E-1   -1.242815E-1   1.461227E-4   3.275149E-6   -3.275149E-6   1.461227E-4   1.461594E-4   1.283995E+0   9.128400E+1   
1.285723E+3   2.041320E+1   2.041320E+1   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   1.063117E-1   -1.260010E-1   1.477900E-4   3.744476E-6   -3.744476E-6   1.477900E-4   1.478374E-4   1.451362E+0   9.145136E+1   
1.307400E+3   2.041781E+1   2.041781E+1   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   1.084206E-1   -1.279878E-1   1.503878E-4   3.483596E-6   -3.483596E-6   1.503878E-4   1.504281E-4   1.326967E+0   9.132697E+1   
1.340545E+3   2.038561E+1   2.038561E+1   4.700000E+1   4.700000E+1   9.000000E+1   4.700000E+1   4.700000E+1   1.083580E-1   -1.271128E-1   1.497792E-4   2.957837E-6   -2.957837E-6   1.497792E-4   1.498084E-4   1.131329E+0   9.113133E+1   
1.361926E+3   2.039431E+1   2.039431E+1   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   1.078104E-1   -1.270994E-1   1.494319E-4   3.354056E-6   -3.354056E-6   1.494319E-4   1.494695E-4   1.285810E+0   9.128581E+1   
1.380971E+3   2.039010E+1   2.039010E+1   4.500000E+1   4.500000E+1   9.000000E+1   4.500000E+1   4.500000E+1   1.080159E-1   -1.273650E-1   1.497320E-4   3.375728E-6   -3.375728E-6   1.497320E-4   1.497700E-4   1.291522E+0   9.129152E+1   
1.403087E+3   2.038821E+1   2.038821E+1   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   1.093474E-1   -1.264680E-1   1.499709E-4   1.804442E-6   -1.804442E-6   1.499709E-4   1.499818E-4   6.893463E-1   9.068935E+1   
1.422162E+3   2.039129E+1   2.039129E+1   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   1.078153E-1   -1.269812E-1   1.493580E-4   3.273199E-6   -3.273199E-6   1.493580E-4   1.493939E-4   1.255443E+0   9.125544E+1   
1.444620E+3   2.036691E+1   2.036691E+1   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   1.096677E-1   -1.260247E-1   1.498802E-4   1.277732E-6   -1.277732E-6   1.498802E-4   1.498857E-4   4.884358E-1   9.048844E+1   
1.463683E+3   2.036230E+1   2.036230E+1   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   1.075938E-1   -1.272650E-1   1.494059E-4   3.622566E-6   -3.622566E-6   1.494059E-4   1.494498E-4   1.388949E+0   9.138895E+1   
1.486082E+3   2.036709E+1   2.036709E+1   3.300000E+1   3.300000E+1   9.000000E+1   3.300000E+1   3.300000E+1   1.084580E-1   -1.264572E-1   1.494141E-4   2.455244E-6   -2.455244E-6   1.494141E-4   1.494343E-4   9.414270E-1   9.094143E+1   
1.507508E+3   2.034179E+1   2.034179E+1   3.100000E+1   3.100000E+1   9.000000E+1   3.100000E+1   3.100000E+1   1.082408E-1   -1.274335E-1   1.499156E-4   3.254126E-6   -3.254126E-6   1.499156E-4   1.499509E-4   1.243489E+0   9.124349E+1   
1.528930E+3   2.035409E+1   2.035409E+1   2.900000E+1   2.900000E+1   9.000000E+1   2.900000E+1   2.900000E+1   1.079632E-1   -1.280427E-1   1.501408E-4   3.857814E-6   -3.857814E-6   1.501408E-4   1.501903E-4   1.471871E+0   9.147187E+1   
1.550361E+3   2.034930E+1   2.034930E+1   2.700000E+1   2.700000E+1   9.000000E+1   2.700000E+1   2.700000E+1   1.080408E-1   -1.275264E-1   1.498525E-4   3.462832E-6   -3.462832E-6   1.498525E-4   1.498925E-4   1.323771E+0   9.132377E+1   
1.571730E+3   2.033071E+1   2.033071E+1   2.500000E+1   2.500000E+1   9.000000E+1   2.500000E+1   2.500000E+1   1.077045E-1   -1.278906E-1   1.498818E-4   3.949621E-6   -3.949621E-6   1.498818E-4   1.499338E-4   1.509485E+0   9.150948E+1   
1.593089E+3   2.033120E+1   2.033120E+1   2.300000E+1   2.300000E+1   9.000000E+1   2.300000E+1   2.300000E+1   1.075959E-1   -1.283302E-1   1.501009E-4   4.317381E-6   -4.317381E-6   1.501009E-4   1.501630E-4   1.647555E+0   9.164755E+1   
1.614528E+3   2.033199E+1   2.033199E+1   2.100000E+1   2.100000E+1   9.000000E+1   2.100000E+1   2.100000E+1   1.084368E-1   -1.276160E-1   1.501557E-4   3.228464E-6   -3.228464E-6   1.501557E-4   1.501904E-4   1.231714E+0   9.123171E+1   
1.635962E+3   2.032809E+1   2.032809E+1   1.900000E+1   1.900000E+1   9.000000E+1   1.900000E+1   1.900000E+1   1.081727E-1   -1.286140E-1   1.506424E-4   4.076307E-6   -4.076307E-6   1.506424E-4   1.506975E-4   1.550017E+0   9.155002E+1   
1.657326E+3   2.032229E+1   2.032229E+1   1.700000E+1   1.700000E+1   9.000000E+1   1.700000E+1   1.700000E+1   1.093038E-1   -1.266398E-1   1.500559E-4   1.948992E-6   -1.948992E-6   1.500559E-4   1.500686E-4   7.441407E-1   9.074414E+1   
1.678661E+3   2.030700E+1   2.030700E+1   1.500000E+1   1.500000E+1   9.000000E+1   1.600000E+1   1.600000E+1   1.081528E-1   -1.287100E-1   1.506925E-4   4.153816E-6   -4.153816E-6   1.506925E-4   1.507498E-4   1.578949E+0   9.157895E+1   
1.700004E+3   2.029510E+1   2.029510E+1   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   1.084675E-1   -1.282811E-1   1.506078E-4   3.640617E-6   -3.640617E-6   1.506078E-4   1.506518E-4   1.384731E+0   9.138473E+1   
1.719108E+3   2.029589E+1   2.029589E+1   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   1.082157E-1   -1.280375E-1   1.502935E-4   3.667657E-6   -3.667657E-6   1.502935E-4   1.503382E-4   1.397929E+0   9.139793E+1   
1.741221E+3   2.029891E+1   2.029891E+1   9.000000E+0   9.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   1.072790E-1   -1.282670E-1   1.498639E-4   4.510440E-6   -4.510440E-6   1.498639E-4   1.499317E-4   1.723906E+0   9.172391E+1   
1.762291E+3   2.029479E+1   2.029479E+1   7.000000E+0   7.000000E+0   9.000000E+1   7.000000E+0   7.000000E+0   1.094367E-1   -1.284520E-1   1.513183E-4   3.035506E-6   -3.035506E-6   1.513183E-4   1.513487E-4   1.149222E+0   9.114922E+1   
1.783368E+3   2.027050E+1   2.027050E+1   5.000000E+0   5.000000E+0   9.000000E+1   6.000000E+0   6.000000E+0   1.093287E-1   -1.287207E-1   1.514266E-4   3.291082E-6   -3.291082E-6   1.514266E-4   1.514623E-4   1.245062E+0   9.124506E+1   
1.804446E+3   2.027169E+1   2.027169E+1   3.000000E+0   3.000000E+0   9.000000E+1   3.000000E+0   3.000000E+0   1.094643E-1   -1.284069E-1   1.513060E-4   2.985617E-6   -2.985617E-6   1.513060E-4   1.513354E-4   1.130432E+0   9.113043E+1   
1.825520E+3   2.025851E+1   2.025851E+1   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   1.097760E-1   -1.288235E-1   1.517701E-4   3.027444E-6   -3.027444E-6   1.517701E-4   1.518002E-4   1.142760E+0   9.114276E+1   
1.844241E+3   2.026049E+1   2.026049E+1   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   1.098229E-1   -1.279464E-1   1.512278E-4   2.419282E-6   -2.419282E-6   1.512278E-4   1.512472E-4   9.165166E-1   9.091652E+1   
1.866230E+3   2.027361E+1   2.027361E+1   -1.000000E+0   -1.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   1.089793E-1   -1.287628E-1   1.512379E-4   3.577022E-6   -3.577022E-6   1.512379E-4   1.512802E-4   1.354886E+0   9.135489E+1   
1.887953E+3   2.024401E+1   2.024401E+1   -3.000000E+0   -3.000000E+0   9.000000E+1   -2.000000E+0   -2.000000E+0   1.088148E-1   -1.300062E-1   1.519461E-4   4.511577E-6   -4.511577E-6   1.519461E-4   1.520130E-4   1.700725E+0   9.170072E+1   
1.909681E+3   2.024182E+1   2.024182E+1   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   1.090311E-1   -1.293073E-1   1.516246E-4   3.894691E-6   -3.894691E-6   1.516246E-4   1.516746E-4   1.471399E+0   9.147140E+1   
1.931723E+3   2.023760E+1   2.023760E+1   -8.000000E+0   -8.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   1.091732E-1   -1.284066E-1   1.511258E-4   3.200751E-6   -3.200751E-6   1.511258E-4   1.511597E-4   1.213308E+0   9.121331E+1   
1.953795E+3   2.024001E+1   2.024001E+1   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   1.099690E-1   -1.285566E-1   1.517155E-4   2.710225E-6   -2.710225E-6   1.517155E-4   1.517397E-4   1.023415E+0   9.102342E+1   
1.976047E+3   2.022549E+1   2.022549E+1   -1.100000E+1   -1.100000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   1.101951E-1   -1.282731E-1   1.516707E-4   2.357666E-6   -2.357666E-6   1.516707E-4   1.516890E-4   8.905703E-1   9.089057E+1   
1.997984E+3   2.020889E+1   2.020889E+1   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   1.082092E-1   -1.284999E-1   1.505906E-4   3.974687E-6   -3.974687E-6   1.505906E-4   1.506430E-4   1.511914E+0   9.151191E+1   
2.020180E+3   2.021301E+1   2.021301E+1   -1.500000E+1   -1.500000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   1.099251E-1   -1.287935E-1   1.518427E-4   2.897493E-6   -2.897493E-6   1.518427E-4   1.518703E-4   1.093197E+0   9.109320E+1   
2.042103E+3   2.021331E+1   2.021331E+1   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   1.099414E-1   -1.292840E-1   1.521722E-4   3.206197E-6   -3.206197E-6   1.521722E-4   1.522060E-4   1.207017E+0   9.120702E+1   
2.064329E+3   2.020510E+1   2.020510E+1   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.800000E+1   -1.800000E+1   1.092741E-1   -1.285416E-1   1.512761E-4   3.214349E-6   -3.214349E-6   1.512761E-4   1.513103E-4   1.217250E+0   9.121725E+1   
2.086610E+3   2.018389E+1   2.018389E+1   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   1.090121E-1   -1.281547E-1   1.508622E-4   3.155203E-6   -3.155203E-6   1.508622E-4   1.508952E-4   1.198136E+0   9.119814E+1   
2.108842E+3   2.018899E+1   2.018899E+1   -2.300000E+1   -2.300000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   1.106727E-1   -1.300513E-1   1.531241E-4   3.166868E-6   -3.166868E-6   1.531241E-4   1.531569E-4   1.184806E+0   9.118481E+1   
2.130756E+3   2.017071E+1   2.017071E+1   -2.500000E+1   -2.500000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   1.096297E-1   -1.294310E-1   1.520752E-4   3.532822E-6   -3.532822E-6   1.520752E-4   1.521162E-4   1.330785E+0   9.133078E+1   
2.152603E+3   2.016839E+1   2.016839E+1   -2.700000E+1   -2.700000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   1.095570E-1   -1.302841E-1   1.525859E-4   4.144367E-6   -4.144367E-6   1.525859E-4   1.526422E-4   1.555821E+0   9.155582E+1   
2.174529E+3   2.016360E+1   2.016360E+1   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   1.099751E-1   -1.294546E-1   1.523042E-4   3.292754E-6   -3.292754E-6   1.523042E-4   1.523398E-4   1.238518E+0   9.123852E+1   
2.196733E+3   2.017031E+1   2.017031E+1   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   1.091235E-1   -1.298289E-1   1.520214E-4   4.167352E-6   -4.167352E-6   1.520214E-4   1.520785E-4   1.570252E+0   9.157025E+1   
2.219008E+3   2.015389E+1   2.015389E+1   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   1.094971E-1   -1.297884E-1   1.522261E-4   3.864491E-6   -3.864491E-6   1.522261E-4   1.522751E-4   1.454229E+0   9.145423E+1   
2.241249E+3   2.014111E+1   2.014111E+1   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   1.109568E-1   -1.286603E-1   1.523938E-4   2.047347E-6   -2.047347E-6   1.523938E-4   1.524076E-4   7.696984E-1   9.076970E+1   
2.263535E+3   2.012759E+1   2.012759E+1   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   1.086719E-1   -1.288382E-1   1.510970E-4   3.853728E-6   -3.853728E-6   1.510970E-4   1.511461E-4   1.461012E+0   9.146101E+1   
2.285801E+3   2.014810E+1   2.014810E+1   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   1.092333E-1   -1.294638E-1   1.518515E-4   3.847439E-6   -3.847439E-6   1.518515E-4   1.519003E-4   1.451384E+0   9.145138E+1   
2.308070E+3   2.012490E+1   2.012490E+1   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   1.099475E-1   -1.300430E-1   1.526703E-4   3.697866E-6   -3.697866E-6   1.526703E-4   1.527151E-4   1.387504E+0   9.138750E+1   
2.330330E+3   2.011730E+1   2.011730E+1   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   1.095735E-1   -1.296853E-1   1.522061E-4   3.740621E-6   -3.740621E-6   1.522061E-4   1.522521E-4   1.407819E+0   9.140782E+1   
2.352598E+3   2.011291E+1   2.011291E+1   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   1.105875E-1   -1.291690E-1   1.524967E-4   2.653112E-6   -2.653112E-6   1.524967E-4   1.525198E-4   9.967216E-1   9.099672E+1   
2.374837E+3   2.011190E+1   2.011190E+1   -4.700000E+1   -4.700000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   1.104408E-1   -1.300700E-1   1.529929E-4   3.350650E-6   -3.350650E-6   1.529929E-4   1.530296E-4   1.254616E+0   9.125462E+1   
2.396751E+3   2.009490E+1   2.009490E+1   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   1.095907E-1   -1.298574E-1   1.523288E-4   3.840428E-6   -3.840428E-6   1.523288E-4   1.523772E-4   1.444203E+0   9.144420E+1   
2.430082E+3   2.010150E+1   2.010150E+1   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   1.114400E-1   -1.315009E-1   1.545426E-4   3.547069E-6   -3.547069E-6   1.545426E-4   1.545833E-4   1.314825E+0   9.131482E+1   
2.451802E+3   2.009701E+1   2.009701E+1   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   1.109311E-1   -1.332337E-1   1.553565E-4   5.056332E-6   -5.056332E-6   1.553565E-4   1.554387E-4   1.864128E+0   9.186413E+1   
2.473509E+3   2.009911E+1   2.009911E+1   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   1.140380E-1   -1.347333E-1   1.582540E-4   3.738781E-6   -3.738781E-6   1.582540E-4   1.582981E-4   1.353372E+0   9.135337E+1   
2.495215E+3   2.010409E+1   2.010409E+1   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   1.136514E-1   -1.358712E-1   1.587561E-4   4.768611E-6   -4.768611E-6   1.587561E-4   1.588277E-4   1.720496E+0   9.172050E+1   
2.517309E+3   2.008529E+1   2.008529E+1   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   1.149749E-1   -1.370759E-1   1.603590E-4   4.577355E-6   -4.577355E-6   1.603590E-4   1.604243E-4   1.635031E+0   9.163503E+1   
2.538982E+3   2.007369E+1   2.007369E+1   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   1.174802E-1   -1.377266E-1   1.623316E-4   3.149796E-6   -3.149796E-6   1.623316E-4   1.623622E-4   1.111597E+0   9.111160E+1   
2.560677E+3   2.006719E+1   2.006719E+1   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   1.166227E-1   -1.412686E-1   1.641083E-4   6.099616E-6   -6.099616E-6   1.641083E-4   1.642216E-4   2.128603E+0   9.212860E+1   
2.582784E+3   2.005969E+1   2.005969E+1   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   1.177541E-1   -1.417493E-1   1.651209E-4   5.577072E-6   -5.577072E-6   1.651209E-4   1.652151E-4   1.934469E+0   9.193447E+1   
2.604455E+3   2.005929E+1   2.005929E+1   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   1.189549E-1   -1.432627E-1   1.668490E-4   5.678343E-6   -5.678343E-6   1.668490E-4   1.669456E-4   1.949185E+0   9.194918E+1   
2.626203E+3   2.006179E+1   2.006179E+1   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   1.199222E-1   -1.450305E-1   1.685983E-4   6.118597E-6   -6.118597E-6   1.685983E-4   1.687093E-4   2.078407E+0   9.207841E+1   
2.647932E+3   2.004760E+1   2.004760E+1   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   1.208610E-1   -1.457987E-1   1.696791E-4   5.926472E-6   -5.926472E-6   1.696791E-4   1.697825E-4   2.000387E+0   9.200039E+1   
2.669665E+3   2.005380E+1   2.005380E+1   -6.510000E+2   -6.510000E+2   9.000000E+1   -6.500000E+2   -6.500000E+2   1.222833E-1   -1.472777E-1   1.715217E-4   5.841468E-6   -5.841468E-6   1.715217E-4   1.716211E-4   1.950553E+0   9.195055E+1   
2.691414E+3   2.004720E+1   2.004720E+1   -7.000000E+2   -7.000000E+2   9.000000E+1   -6.990000E+2   -6.990000E+2   1.226334E-1   -1.493394E-1   1.730808E-4   6.930402E-6   -6.930402E-6   1.730808E-4   1.732195E-4   2.292979E+0   9.229298E+1   
2.713138E+3   2.005279E+1   2.005279E+1   -7.500000E+2   -7.500000E+2   9.000000E+1   -7.490000E+2   -7.490000E+2   1.232509E-1   -1.508696E-1   1.744593E-4   7.474075E-6   -7.474075E-6   1.744593E-4   1.746193E-4   2.453130E+0   9.245313E+1   
2.734870E+3   2.002361E+1   2.002361E+1   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   1.244253E-1   -1.528776E-1   1.764931E-4   7.918196E-6   -7.918196E-6   1.764931E-4   1.766707E-4   2.568798E+0   9.256880E+1   
2.756557E+3   2.002590E+1   2.002590E+1   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   1.260403E-1   -1.538983E-1   1.781564E-4   7.391032E-6   -7.391032E-6   1.781564E-4   1.783096E-4   2.375623E+0   9.237562E+1   
2.778192E+3   2.002090E+1   2.002090E+1   -9.000000E+2   -9.000000E+2   9.000000E+1   -8.990000E+2   -8.990000E+2   1.264968E-1   -1.542088E-1   1.786408E-4   7.256365E-6   -7.256365E-6   1.786408E-4   1.787881E-4   2.326068E+0   9.232607E+1   
2.799879E+3   2.001150E+1   2.001150E+1   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   1.284241E-1   -1.561615E-1   1.811041E-4   7.107546E-6   -7.107546E-6   1.811041E-4   1.812435E-4   2.247456E+0   9.224746E+1   
2.821509E+3   1.999969E+1   1.999969E+1   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   1.284321E-1   -1.584296E-1   1.825862E-4   8.584469E-6   -8.584469E-6   1.825862E-4   1.827879E-4   2.691834E+0   9.269183E+1   
2.844044E+3   2.000280E+1   2.000280E+1   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   1.298979E-1   -1.585646E-1   1.835804E-4   7.588527E-6   -7.588527E-6   1.835804E-4   1.837372E-4   2.367046E+0   9.236705E+1   
2.865911E+3   2.000009E+1   2.000009E+1   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   1.305640E-1   -1.604965E-1   1.852504E-4   8.358913E-6   -8.358913E-6   1.852504E-4   1.854389E-4   2.583561E+0   9.258356E+1   
2.887782E+3   1.999609E+1   1.999609E+1   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   1.301255E-1   -1.626864E-1   1.864056E-4   1.011486E-5   -1.011486E-5   1.864056E-4   1.866798E-4   3.105974E+0   9.310597E+1   
2.910147E+3   1.997131E+1   1.997131E+1   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   1.323869E-1   -1.635613E-1   1.883735E-4   9.014305E-6   -9.014305E-6   1.883735E-4   1.885891E-4   2.739705E+0   9.273970E+1   
2.932192E+3   1.997341E+1   1.997341E+1   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   1.323529E-1   -1.654291E-1   1.895689E-4   1.026056E-5   -1.026056E-5   1.895689E-4   1.898464E-4   3.098154E+0   9.309815E+1   
2.954293E+3   1.997939E+1   1.997939E+1   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   1.338071E-1   -1.662559E-1   1.910065E-4   9.725551E-6   -9.725551E-6   1.910065E-4   1.912539E-4   2.914834E+0   9.291483E+1   
2.976618E+3   1.998071E+1   1.998071E+1   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   1.361970E-1   -1.679071E-1   1.935594E-4   9.037375E-6   -9.037375E-6   1.935594E-4   1.937703E-4   2.673224E+0   9.267322E+1   
2.998741E+3   1.996191E+1   1.996191E+1   -1.399000E+3   -1.399000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   1.357202E-1   -1.692772E-1   1.941571E-4   1.028574E-5   -1.028574E-5   1.941571E-4   1.944293E-4   3.032490E+0   9.303249E+1   
3.020876E+3   1.995120E+1   1.995120E+1   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   1.378377E-1   -1.699187E-1   1.958840E-4   9.139000E-6   -9.139000E-6   1.958840E-4   1.960970E-4   2.671208E+0   9.267121E+1   
3.044016E+3   1.996121E+1   1.996121E+1   -1.499000E+3   -1.499000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   1.369235E-1   -1.719727E-1   1.966565E-4   1.115802E-5   -1.115802E-5   1.966565E-4   1.969728E-4   3.247403E+0   9.324740E+1   
3.066093E+3   1.993990E+1   1.993990E+1   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.548000E+3   -1.548000E+3   1.382629E-1   -1.732281E-1   1.983022E-4   1.098807E-5   -1.098807E-5   1.983022E-4   1.986064E-4   3.171558E+0   9.317156E+1   
3.088687E+3   1.994161E+1   1.994161E+1   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   1.390164E-1   -1.755612E-1   2.002876E-4   1.195612E-5   -1.195612E-5   2.002876E-4   2.006442E-4   3.416204E+0   9.341620E+1   
3.111772E+3   1.992281E+1   1.992281E+1   -1.650000E+3   -1.650000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   1.398954E-1   -1.762221E-1   2.012614E-4   1.173805E-5   -1.173805E-5   2.012614E-4   2.016034E-4   3.337848E+0   9.333785E+1   
3.133797E+3   1.992458E+1   1.992458E+1   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.698000E+3   -1.698000E+3   1.408363E-1   -1.786378E-1   2.034165E-4   1.262141E-5   -1.262141E-5   2.034165E-4   2.038076E-4   3.550488E+0   9.355049E+1   
3.155912E+3   1.991299E+1   1.991299E+1   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.748000E+3   -1.748000E+3   1.402534E-1   -1.805402E-1   2.042951E-4   1.429630E-5   -1.429630E-5   2.042951E-4   2.047947E-4   4.002956E+0   9.400296E+1   
3.179547E+3   1.991131E+1   1.991131E+1   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.799000E+3   -1.799000E+3   1.426642E-1   -1.811099E-1   2.061566E-4   1.288567E-5   -1.288567E-5   2.061566E-4   2.065589E-4   3.576578E+0   9.357658E+1   
3.201676E+3   1.990389E+1   1.990389E+1   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.848000E+3   -1.848000E+3   1.427212E-1   -1.836219E-1   2.078279E-4   1.448575E-5   -1.448575E-5   2.078279E-4   2.083321E-4   3.987108E+0   9.398711E+1   
3.224067E+3   1.990130E+1   1.990130E+1   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   1.449998E-1   -1.843156E-1   2.096884E-4   1.325396E-5   -1.325396E-5   2.096884E-4   2.101069E-4   3.616732E+0   9.361673E+1   
3.247397E+3   1.989260E+1   1.989260E+1   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.948000E+3   -1.948000E+3   1.436996E-1   -1.855382E-1   2.096809E-4   1.501497E-5   -1.501497E-5   2.096809E-4   2.102178E-4   4.095883E+0   9.409588E+1   
3.269787E+3   1.988339E+1   1.988339E+1   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   1.457523E-1   -1.870048E-1   2.119051E-4   1.445548E-5   -1.445548E-5   2.119051E-4   2.123976E-4   3.902485E+0   9.390249E+1   
3.307330E+3   1.986749E+1   1.986749E+1   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.556320E-1   -2.025281E-1   2.281234E-4   1.729690E-5   -1.729690E-5   2.281234E-4   2.287782E-4   4.336016E+0   9.433602E+1   
3.333431E+3   1.986810E+1   1.986810E+1   -2.999000E+3   -2.999000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.643759E-1   -2.181491E-1   2.437030E-4   2.104218E-5   -2.104218E-5   2.437030E-4   2.446098E-4   4.934882E+0   9.493488E+1   
3.359139E+3   1.987289E+1   1.987289E+1   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.749688E-1   -2.353727E-1   2.614696E-4   2.446766E-5   -2.446766E-5   2.614696E-4   2.626120E-4   5.346024E+0   9.534602E+1   
3.384738E+3   1.984130E+1   1.984130E+1   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   1.855349E-1   -2.533956E-1   2.797402E-4   2.843556E-5   -2.843556E-5   2.797402E-4   2.811818E-4   5.804172E+0   9.580417E+1   
3.410969E+3   1.986199E+1   1.986199E+1   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   1.976130E-1   -2.689015E-1   2.973063E-4   2.963953E-5   -2.963953E-5   2.973063E-4   2.987801E-4   5.693210E+0   9.569321E+1   
3.436111E+3   1.985790E+1   1.985790E+1   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   2.049159E-1   -2.827067E-1   3.108125E-4   3.326354E-5   -3.326354E-5   3.108125E-4   3.125873E-4   6.108615E+0   9.610862E+1   
3.461380E+3   1.985500E+1   1.985500E+1   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   2.108560E-1   -2.953051E-1   3.226901E-4   3.710652E-5   -3.710652E-5   3.226901E-4   3.248166E-4   6.559698E+0   9.655970E+1   
3.487596E+3   1.984429E+1   1.984429E+1   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   2.162414E-1   -3.042262E-1   3.318299E-4   3.895564E-5   -3.895564E-5   3.318299E-4   3.341087E-4   6.695673E+0   9.669567E+1   
3.512805E+3   1.984060E+1   1.984060E+1   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   2.138825E-1   -3.059349E-1   3.314843E-4   4.181744E-5   -4.181744E-5   3.314843E-4   3.341116E-4   7.190002E+0   9.719000E+1   
3.537497E+3   1.982861E+1   1.982861E+1   -7.000000E+3   -7.000000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.968003E-1   -2.867317E-1   3.084164E-4   4.189746E-5   -4.189746E-5   3.084164E-4   3.112492E-4   7.736106E+0   9.773611E+1   
3.562665E+3   1.982031E+1   1.982031E+1   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.807276E-1   -2.674200E-1   2.859021E-4   4.115985E-5   -4.115985E-5   2.859021E-4   2.888497E-4   8.192291E+0   9.819229E+1   
3.587874E+3   1.980639E+1   1.980639E+1   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.643568E-1   -2.511821E-1   2.652053E-4   4.265231E-5   -4.265231E-5   2.652053E-4   2.686132E-4   9.136501E+0   9.913650E+1   
3.613542E+3   1.979061E+1   1.979061E+1   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.564428E-1   -2.420890E-1   2.543903E-4   4.256099E-5   -4.256099E-5   2.543903E-4   2.579261E-4   9.497953E+0   9.949795E+1   
3.639283E+3   1.980190E+1   1.980190E+1   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.528113E-1   -2.415739E-1   2.518096E-4   4.491017E-5   -4.491017E-5   2.518096E-4   2.557831E-4   1.011236E+1   1.001124E+2   
3.664530E+3   1.979791E+1   1.979791E+1   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.474385E-1   -2.395969E-1   2.472003E-4   4.759162E-5   -4.759162E-5   2.472003E-4   2.517398E-4   1.089740E+1   1.008974E+2   
3.689690E+3   1.979699E+1   1.979699E+1   -9.999000E+3   -9.999000E+3   9.000000E+1   -9.998000E+3   -9.998000E+3   1.613377E-1   -2.542226E-1   2.653190E-4   4.687320E-5   -4.687320E-5   2.653190E-4   2.694277E-4   1.001891E+1   1.000189E+2   
3.726271E+3   1.978909E+1   1.978909E+1   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.384918E-1   -2.243395E-1   2.317320E-4   4.423399E-5   -4.423399E-5   2.317320E-4   2.359161E-4   1.080686E+1   1.008069E+2   
3.750452E+3   1.978271E+1   1.978271E+1   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.218112E-1   -2.044412E-1   2.084598E-4   4.356259E-5   -4.356259E-5   2.084598E-4   2.129628E-4   1.180344E+1   1.018034E+2   
3.774604E+3   1.977810E+1   1.977810E+1   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.091867E-1   -1.873353E-1   1.895138E-4   4.171667E-5   -4.171667E-5   1.895138E-4   1.940509E-4   1.241424E+1   1.024142E+2   
3.798836E+3   1.978011E+1   1.978011E+1   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   9.318230E-2   -1.670667E-1   1.664185E-4   4.030300E-5   -4.030300E-5   1.664185E-4   1.712292E-4   1.361370E+1   1.036137E+2   
3.823524E+3   1.976809E+1   1.976809E+1   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   8.141729E-2   -1.491461E-1   1.474732E-4   3.728874E-5   -3.728874E-5   1.474732E-4   1.521145E-4   1.418988E+1   1.041899E+2   
3.848712E+3   1.976751E+1   1.976751E+1   -7.000000E+3   -7.000000E+3   9.000000E+1   -6.999000E+3   -6.999000E+3   7.046140E-2   -1.325483E-1   1.298898E-4   3.454089E-5   -3.454089E-5   1.298898E-4   1.344040E-4   1.489171E+1   1.048917E+2   
3.873355E+3   1.976449E+1   1.976449E+1   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   5.695793E-2   -1.143487E-1   1.096882E-4   3.263013E-5   -3.263013E-5   1.096882E-4   1.144387E-4   1.656673E+1   1.065667E+2   
3.897562E+3   1.976440E+1   1.976440E+1   -5.999000E+3   -5.999000E+3   9.000000E+1   -5.998000E+3   -5.998000E+3   4.906471E-2   -9.958801E-2   9.519471E-5   2.881804E-5   -2.881804E-5   9.519471E-5   9.946111E-5   1.684250E+1   1.068425E+2   
3.922332E+3   1.976461E+1   1.976461E+1   -5.499000E+3   -5.499000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   4.159483E-2   -8.585628E-2   8.163315E-5   2.536558E-5   -2.536558E-5   8.163315E-5   8.548324E-5   1.726140E+1   1.072614E+2   
3.947115E+3   1.976241E+1   1.976241E+1   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   3.061839E-2   -6.973586E-2   6.434794E-5   2.294502E-5   -2.294502E-5   6.434794E-5   6.831641E-5   1.962509E+1   1.096251E+2   
3.971298E+3   1.977389E+1   1.977389E+1   -4.499000E+3   -4.499000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   1.549709E-2   -4.898711E-2   4.148581E-5   2.056426E-5   -2.056426E-5   4.148581E-5   4.630293E-5   2.636733E+1   1.163673E+2   
3.996020E+3   1.976711E+1   1.976711E+1   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   7.204757E-3   -3.525647E-2   2.741648E-5   1.772082E-5   -1.772082E-5   2.741648E-5   3.264492E-5   3.287687E+1   1.228769E+2   
4.020702E+3   1.977068E+1   1.977068E+1   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   -1.605455E-3   -1.886906E-2   1.129665E-5   1.352351E-5   -1.352351E-5   1.129665E-5   1.762100E-5   5.012682E+1   1.401268E+2   
4.044857E+3   1.976940E+1   1.976940E+1   -2.999000E+3   -2.999000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   -1.325045E-2   -3.481193E-3   -5.924783E-6   1.207635E-5   -1.207635E-5   -5.924783E-6   1.345144E-5   1.161331E+2   2.061331E+2   
4.069511E+3   1.977542E+1   1.977542E+1   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   -2.092674E-2   1.150202E-2   -2.042904E-5   7.958367E-6   -7.958367E-6   -2.042904E-5   2.192444E-5   1.587160E+2   2.487160E+2   
4.093690E+3   1.977709E+1   1.977709E+1   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   -3.222629E-2   2.910529E-2   -3.887976E-5   4.807348E-6   -4.807348E-6   -3.887976E-5   3.917584E-5   1.729514E+2   2.629514E+2   
4.127373E+3   1.979101E+1   1.979101E+1   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.948000E+3   -1.948000E+3   -3.338965E-2   3.123412E-2   -4.098550E-5   4.276038E-6   -4.276038E-6   -4.098550E-5   4.120795E-5   1.740439E+2   2.640439E+2   
4.149425E+3   1.977661E+1   1.977661E+1   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   -3.317427E-2   3.301566E-2   -4.201264E-5   2.952015E-6   -2.952015E-6   -4.201264E-5   4.211622E-5   1.759807E+2   2.659807E+2   
4.171528E+3   1.978521E+1   1.978521E+1   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.848000E+3   -1.848000E+3   -3.453705E-2   3.555191E-2   -4.450700E-5   2.301838E-6   -2.301838E-6   -4.450700E-5   4.456649E-5   1.770394E+2   2.670394E+2   
4.193300E+3   1.979269E+1   1.979269E+1   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.798000E+3   -1.798000E+3   -3.439410E-2   3.768842E-2   -4.581011E-5   7.993193E-7   -7.993193E-7   -4.581011E-5   4.581708E-5   1.790004E+2   2.690004E+2   
4.215394E+3   1.977889E+1   1.977889E+1   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   -3.624373E-2   3.829894E-2   -4.735126E-5   1.768228E-6   -1.768228E-6   -4.735126E-5   4.738426E-5   1.778614E+2   2.678614E+2   
4.237399E+3   1.979171E+1   1.979171E+1   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   -3.688831E-2   3.984025E-2   -4.875361E-5   1.237315E-6   -1.237315E-6   -4.875361E-5   4.876931E-5   1.785462E+2   2.685462E+2   
4.259180E+3   1.978719E+1   1.978719E+1   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   -3.735249E-2   3.983874E-2   -4.903960E-5   1.581616E-6   -1.581616E-6   -4.903960E-5   4.906510E-5   1.781527E+2   2.681527E+2   
4.281016E+3   1.979199E+1   1.979199E+1   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.599000E+3   -1.599000E+3   -3.831735E-2   4.169483E-2   -5.084498E-5   1.081801E-6   -1.081801E-6   -5.084498E-5   5.085649E-5   1.787811E+2   2.687811E+2   
4.303179E+3   1.978781E+1   1.978781E+1   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   -3.854161E-2   4.420501E-2   -5.261848E-5   -3.934139E-7   3.934139E-7   -5.261848E-5   5.261995E-5   -1.795716E+2   -8.957162E+1   
4.325048E+3   1.978359E+1   1.978359E+1   -1.499000E+3   -1.499000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   -3.984825E-2   4.532204E-2   -5.415382E-5   -1.572682E-7   1.572682E-7   -5.415382E-5   5.415405E-5   -1.798336E+2   -8.983361E+1   
4.347129E+3   1.978951E+1   1.978951E+1   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   -4.155616E-2   4.715001E-2   -5.640027E-5   -8.911695E-8   8.911695E-8   -5.640027E-5   5.640034E-5   -1.799095E+2   -8.990947E+1   
4.369142E+3   1.978399E+1   1.978399E+1   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   -4.207218E-2   4.670637E-2   -5.643035E-5   5.825874E-7   -5.825874E-7   -5.643035E-5   5.643336E-5   1.794085E+2   2.694085E+2   
4.391013E+3   1.979571E+1   1.979571E+1   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   -4.328219E-2   4.929792E-2   -5.886629E-5   -2.167393E-7   2.167393E-7   -5.886629E-5   5.886668E-5   -1.797890E+2   -8.978904E+1   
4.413119E+3   1.979571E+1   1.979571E+1   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   -4.427314E-2   4.948811E-2   -5.960281E-5   3.918650E-7   -3.918650E-7   -5.960281E-5   5.960410E-5   1.796233E+2   2.696233E+2   
4.435182E+3   1.979061E+1   1.979061E+1   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   -4.508736E-2   5.371237E-2   -6.285741E-5   -1.767614E-6   1.767614E-6   -6.285741E-5   6.288226E-5   -1.783892E+2   -8.838921E+1   
4.457017E+3   1.979180E+1   1.979180E+1   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   -4.547426E-2   5.473828E-2   -6.376477E-5   -2.152165E-6   2.152165E-6   -6.376477E-5   6.380108E-5   -1.780669E+2   -8.806691E+1   
4.479140E+3   1.978051E+1   1.978051E+1   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   -4.580990E-2   5.597589E-2   -6.477833E-5   -2.713030E-6   2.713030E-6   -6.477833E-5   6.483511E-5   -1.776018E+2   -8.760175E+1   
4.501121E+3   1.979131E+1   1.979131E+1   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.100000E+3   -1.100000E+3   -4.716227E-2   5.630692E-2   -6.583002E-5   -1.929197E-6   1.929197E-6   -6.583002E-5   6.585828E-5   -1.783214E+2   -8.832139E+1   
4.522940E+3   1.978301E+1   1.978301E+1   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   -4.826706E-2   5.798751E-2   -6.760761E-5   -2.210781E-6   2.210781E-6   -6.760761E-5   6.764374E-5   -1.781271E+2   -8.812708E+1   
4.544962E+3   1.978130E+1   1.978130E+1   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   -4.931324E-2   5.918432E-2   -6.903387E-5   -2.219434E-6   2.219434E-6   -6.903387E-5   6.906954E-5   -1.781586E+2   -8.815858E+1   
4.566840E+3   1.978430E+1   1.978430E+1   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   -4.988390E-2   6.095636E-2   -7.054079E-5   -2.955861E-6   2.955861E-6   -7.054079E-5   7.060269E-5   -1.776005E+2   -8.760055E+1   
4.588509E+3   1.978381E+1   1.978381E+1   -9.000000E+2   -9.000000E+2   9.000000E+1   -8.990000E+2   -8.990000E+2   -5.124206E-2   6.278147E-2   -7.256915E-5   -3.144532E-6   3.144532E-6   -7.256915E-5   7.263724E-5   -1.775188E+2   -8.751884E+1   
4.610433E+3   1.977831E+1   1.977831E+1   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   -5.205385E-2   6.403931E-2   -7.389025E-5   -3.366447E-6   3.366447E-6   -7.389025E-5   7.396689E-5   -1.773914E+2   -8.739140E+1   
4.632061E+3   1.976309E+1   1.976309E+1   -8.000000E+2   -8.000000E+2   9.000000E+1   -8.000000E+2   -8.000000E+2   -5.266898E-2   6.561744E-2   -7.529837E-5   -3.943218E-6   3.943218E-6   -7.529837E-5   7.540155E-5   -1.770023E+2   -8.700228E+1   
4.653702E+3   1.976910E+1   1.976910E+1   -7.500000E+2   -7.500000E+2   9.000000E+1   -7.490000E+2   -7.490000E+2   -5.427442E-2   6.696028E-2   -7.716551E-5   -3.633697E-6   3.633697E-6   -7.716551E-5   7.725102E-5   -1.773040E+2   -8.730395E+1   
4.675633E+3   1.976681E+1   1.976681E+1   -7.000000E+2   -7.000000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   -5.531170E-2   6.834882E-2   -7.871114E-5   -3.774278E-6   3.774278E-6   -7.871114E-5   7.880158E-5   -1.772547E+2   -8.725471E+1   
4.697563E+3   1.976541E+1   1.976541E+1   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.490000E+2   -6.490000E+2   -5.592406E-2   7.109983E-2   -8.088144E-5   -5.119891E-6   5.119891E-6   -8.088144E-5   8.104332E-5   -1.763779E+2   -8.637794E+1   
4.719246E+3   1.976760E+1   1.976760E+1   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   -5.737272E-2   7.195210E-2   -8.233214E-5   -4.605604E-6   4.605604E-6   -8.233214E-5   8.246086E-5   -1.767983E+2   -8.679825E+1   
4.740882E+3   1.977361E+1   1.977361E+1   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.500000E+2   -5.500000E+2   -5.784793E-2   7.328113E-2   -8.349152E-5   -5.123008E-6   5.123008E-6   -8.349152E-5   8.364855E-5   -1.764888E+2   -8.648875E+1   
4.762502E+3   1.977169E+1   1.977169E+1   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   -5.835322E-2   7.465097E-2   -8.469608E-5   -5.644840E-6   5.644840E-6   -8.469608E-5   8.488398E-5   -1.761870E+2   -8.618698E+1   
4.784183E+3   1.979141E+1   1.979141E+1   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   -5.922482E-2   7.562379E-2   -8.586853E-5   -5.636182E-6   5.636182E-6   -8.586853E-5   8.605330E-5   -1.762446E+2   -8.624464E+1   
4.805814E+3   1.977050E+1   1.977050E+1   -3.990000E+2   -3.990000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   -6.061091E-2   7.714151E-2   -8.771395E-5   -5.603228E-6   5.603228E-6   -8.771395E-5   8.789273E-5   -1.763449E+2   -8.634487E+1   
4.827550E+3   1.977801E+1   1.977801E+1   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   -6.103736E-2   7.787476E-2   -8.845515E-5   -5.767189E-6   5.767189E-6   -8.845515E-5   8.864296E-5   -1.762697E+2   -8.626965E+1   
4.849281E+3   1.975948E+1   1.975948E+1   -2.990000E+2   -2.990000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   -6.202155E-2   7.963634E-2   -9.021093E-5   -6.190926E-6   6.190926E-6   -9.021093E-5   9.042311E-5   -1.760741E+2   -8.607410E+1   
4.870906E+3   1.977999E+1   1.977999E+1   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   -6.221819E-2   8.315709E-2   -9.262553E-5   -8.347250E-6   8.347250E-6   -9.262553E-5   9.300089E-5   -1.748505E+2   -8.485052E+1   
4.892586E+3   1.978481E+1   1.978481E+1   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   -6.329904E-2   8.294326E-2   -9.315449E-5   -7.408024E-6   7.408024E-6   -9.315449E-5   9.344859E-5   -1.754532E+2   -8.545318E+1   
4.914227E+3   1.977249E+1   1.977249E+1   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   -6.375982E-2   8.413391E-2   -9.421483E-5   -7.845626E-6   7.845626E-6   -9.421483E-5   9.454093E-5   -1.752397E+2   -8.523975E+1   
4.935903E+3   1.978820E+1   1.978820E+1   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   -6.419211E-2   8.588601E-2   -9.562321E-5   -8.671370E-6   8.671370E-6   -9.562321E-5   9.601558E-5   -1.748184E+2   -8.481844E+1   
4.957383E+3   1.977639E+1   1.977639E+1   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   -6.622890E-2   8.730861E-2   -9.780898E-5   -8.094955E-6   8.094955E-6   -9.780898E-5   9.814339E-5   -1.752688E+2   -8.526882E+1   
4.990373E+3   1.976919E+1   1.976919E+1   -4.700000E+1   -4.700000E+1   9.000000E+1   -4.600000E+1   -4.600000E+1   -6.503302E-2   8.739820E-2   -9.712798E-5   -9.038030E-6   9.038030E-6   -9.712798E-5   9.754758E-5   -1.746838E+2   -8.468378E+1   
5.011642E+3   1.976119E+1   1.976119E+1   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   -6.659829E-2   8.644009E-2   -9.747169E-5   -7.253927E-6   7.253927E-6   -9.747169E-5   9.774124E-5   -1.757438E+2   -8.574384E+1   
5.033851E+3   1.975631E+1   1.975631E+1   -4.300000E+1   -4.300000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   -6.751651E-2   8.654745E-2   -9.810930E-5   -6.644967E-6   6.644967E-6   -9.810930E-5   9.833407E-5   -1.761253E+2   -8.612526E+1   
5.055134E+3   1.974041E+1   1.974041E+1   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   -6.601477E-2   8.744942E-2   -9.776830E-5   -8.345392E-6   8.345392E-6   -9.776830E-5   9.812383E-5   -1.751211E+2   -8.512112E+1   
5.077305E+3   1.975640E+1   1.975640E+1   -3.900000E+1   -3.900000E+1   9.000000E+1   -3.800000E+1   -3.800000E+1   -6.593254E-2   8.710827E-2   -9.749527E-5   -8.183172E-6   8.183172E-6   -9.749527E-5   9.783809E-5   -1.752022E+2   -8.520218E+1   
5.098545E+3   1.975219E+1   1.975219E+1   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   -6.591198E-2   8.664594E-2   -9.718145E-5   -7.896125E-6   7.896125E-6   -9.718145E-5   9.750171E-5   -1.753548E+2   -8.535484E+1   
5.120780E+3   1.976879E+1   1.976879E+1   -3.500000E+1   -3.500000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   -6.619240E-2   8.741844E-2   -9.785795E-5   -8.193753E-6   8.193753E-6   -9.785795E-5   9.820038E-5   -1.752137E+2   -8.521373E+1   
5.142054E+3   1.975430E+1   1.975430E+1   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   -6.664981E-2   8.725492E-2   -9.803423E-5   -7.748532E-6   7.748532E-6   -9.803423E-5   9.833997E-5   -1.754808E+2   -8.548079E+1   
5.164289E+3   1.975430E+1   1.975430E+1   -3.100000E+1   -3.100000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   -6.672530E-2   8.694935E-2   -9.788189E-5   -7.492923E-6   7.492923E-6   -9.788189E-5   9.816827E-5   -1.756225E+2   -8.562251E+1   
5.185553E+3   1.976019E+1   1.976019E+1   -2.900000E+1   -2.900000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   -6.706645E-2   8.763965E-2   -9.854239E-5   -7.691904E-6   7.691904E-6   -9.854239E-5   9.884214E-5   -1.755367E+2   -8.553672E+1   
5.206752E+3   1.974111E+1   1.974111E+1   -2.700000E+1   -2.700000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   -6.654705E-2   8.745250E-2   -9.809938E-5   -7.953712E-6   7.953712E-6   -9.809938E-5   9.842129E-5   -1.753647E+2   -8.536471E+1   
5.227919E+3   1.974941E+1   1.974941E+1   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   -6.613749E-2   8.740402E-2   -9.781460E-5   -8.224938E-6   8.224938E-6   -9.781460E-5   9.815979E-5   -1.751935E+2   -8.519348E+1   
5.250148E+3   1.974600E+1   1.974600E+1   -2.300000E+1   -2.300000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   -6.622278E-2   8.763227E-2   -9.801599E-5   -8.311083E-6   8.311083E-6   -9.801599E-5   9.836772E-5   -1.751533E+2   -8.515330E+1   
5.271432E+3   1.973989E+1   1.973989E+1   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   -6.713609E-2   8.725459E-2   -9.833466E-5   -7.388648E-6   7.388648E-6   -9.833466E-5   9.861185E-5   -1.757030E+2   -8.570300E+1   
5.293705E+3   1.973589E+1   1.973589E+1   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   -6.710725E-2   8.743256E-2   -9.843274E-5   -7.526327E-6   7.526327E-6   -9.843274E-5   9.872006E-5   -1.756276E+2   -8.562758E+1   
5.315948E+3   1.973550E+1   1.973550E+1   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   -6.776134E-2   8.806364E-2   -9.924814E-5   -7.455131E-6   7.455131E-6   -9.924814E-5   9.952775E-5   -1.757042E+2   -8.570423E+1   
5.338138E+3   1.974081E+1   1.974081E+1   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   -6.796933E-2   8.749544E-2   -9.900667E-5   -6.929822E-6   6.929822E-6   -9.900667E-5   9.924890E-5   -1.759962E+2   -8.599620E+1   
5.360414E+3   1.974719E+1   1.974719E+1   -1.300000E+1   -1.300000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   -6.729132E-2   8.801239E-2   -9.892418E-5   -7.769259E-6   7.769259E-6   -9.892418E-5   9.922880E-5   -1.755093E+2   -8.550935E+1   
5.381683E+3   1.974249E+1   1.974249E+1   -1.100000E+1   -1.100000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   -6.748552E-2   8.860451E-2   -9.942988E-5   -8.012742E-6   8.012742E-6   -9.942988E-5   9.975222E-5   -1.753927E+2   -8.539267E+1   
5.402786E+3   1.975210E+1   1.975210E+1   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   -6.693268E-2   8.812345E-2   -9.877478E-5   -8.107134E-6   8.107134E-6   -9.877478E-5   9.910692E-5   -1.753079E+2   -8.530785E+1   
5.424911E+3   1.973708E+1   1.973708E+1   -8.000000E+0   -8.000000E+0   9.000000E+1   -6.000000E+0   -6.000000E+0   -6.689250E-2   8.813605E-2   -9.875815E-5   -8.145087E-6   8.145087E-6   -9.875815E-5   9.909346E-5   -1.752852E+2   -8.528520E+1   
5.446999E+3   1.974520E+1   1.974520E+1   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   -6.645409E-2   8.857076E-2   -9.877022E-5   -8.753550E-6   8.753550E-6   -9.877022E-5   9.915735E-5   -1.749354E+2   -8.493537E+1   
5.469039E+3   1.973239E+1   1.973239E+1   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   -6.541466E-2   8.795288E-2   -9.772518E-5   -9.118393E-6   9.118393E-6   -9.772518E-5   9.814966E-5   -1.746694E+2   -8.466937E+1   
5.491176E+3   1.973309E+1   1.973309E+1   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   -6.708792E-2   8.898310E-2   -9.943064E-5   -8.554322E-6   8.554322E-6   -9.943064E-5   9.979794E-5   -1.750828E+2   -8.508278E+1   
5.513205E+3   1.972360E+1   1.972360E+1   0.000000E+0   0.000000E+0   9.000000E+1   0.000000E+0   0.000000E+0   -6.694555E-2   8.804154E-2   -9.872940E-5   -8.044062E-6   8.044062E-6   -9.872940E-5   9.905655E-5   -1.753421E+2   -8.534207E+1   
5.535232E+3   1.971649E+1   1.971649E+1   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   -6.719468E-2   8.796361E-2   -9.883266E-5   -7.808852E-6   7.808852E-6   -9.883266E-5   9.914067E-5   -1.754824E+2   -8.548240E+1   
5.556714E+3   1.972030E+1   1.972030E+1   3.000000E+0   3.000000E+0   9.000000E+1   4.000000E+0   4.000000E+0   -6.720143E-2   8.724878E-2   -9.837127E-5   -7.336522E-6   7.336522E-6   -9.837127E-5   9.864447E-5   -1.757348E+2   -8.573478E+1   
5.578441E+3   1.972021E+1   1.972021E+1   5.000000E+0   5.000000E+0   9.000000E+1   6.000000E+0   6.000000E+0   -6.736587E-2   8.799767E-2   -9.896068E-5   -7.704500E-6   7.704500E-6   -9.896068E-5   9.926014E-5   -1.755483E+2   -8.554827E+1   
5.600156E+3   1.971230E+1   1.971230E+1   7.000000E+0   7.000000E+0   9.000000E+1   8.000000E+0   8.000000E+0   -6.715788E-2   8.805075E-2   -9.886666E-5   -7.893037E-6   7.893037E-6   -9.886666E-5   9.918123E-5   -1.754355E+2   -8.543546E+1   
5.621903E+3   1.970211E+1   1.970211E+1   9.000000E+0   9.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   -6.716859E-2   8.822011E-2   -9.898359E-5   -7.995838E-6   7.995838E-6   -9.898359E-5   9.930601E-5   -1.753817E+2   -8.538171E+1   
5.643936E+3   1.970571E+1   1.970571E+1   1.100000E+1   1.100000E+1   9.000000E+1   1.100000E+1   1.100000E+1   -6.724192E-2   8.841737E-2   -9.915740E-5   -8.070564E-6   8.070564E-6   -9.915740E-5   9.948529E-5   -1.753469E+2   -8.534687E+1   
5.665978E+3   1.969390E+1   1.969390E+1   1.300000E+1   1.300000E+1   9.000000E+1   1.300000E+1   1.300000E+1   -6.789081E-2   8.870881E-2   -9.974838E-5   -7.781168E-6   7.781168E-6   -9.974838E-5   1.000514E-4   -1.755395E+2   -8.553951E+1   
5.688082E+3   1.969470E+1   1.969470E+1   1.500000E+1   1.500000E+1   9.000000E+1   1.600000E+1   1.600000E+1   -6.790613E-2   8.827930E-2   -9.947812E-5   -7.489028E-6   7.489028E-6   -9.947812E-5   9.975962E-5   -1.756947E+2   -8.569471E+1   
5.710078E+3   1.969201E+1   1.969201E+1   1.700000E+1   1.700000E+1   9.000000E+1   1.700000E+1   1.700000E+1   -6.784355E-2   8.840969E-2   -9.952435E-5   -7.620558E-6   7.620558E-6   -9.952435E-5   9.981567E-5   -1.756214E+2   -8.562142E+1   
5.732138E+3   1.968710E+1   1.968710E+1   1.900000E+1   1.900000E+1   9.000000E+1   1.900000E+1   1.900000E+1   -6.734196E-2   8.921840E-2   -9.974095E-5   -8.520263E-6   8.520263E-6   -9.974095E-5   1.001042E-4   -1.751174E+2   -8.511742E+1   
5.754221E+3   1.967440E+1   1.967440E+1   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   -6.789724E-2   8.857597E-2   -9.966584E-5   -7.689557E-6   7.689557E-6   -9.966584E-5   9.996204E-5   -1.755882E+2   -8.558818E+1   
5.776050E+3   1.967809E+1   1.967809E+1   2.300000E+1   2.300000E+1   9.000000E+1   2.400000E+1   2.400000E+1   -6.813839E-2   8.818052E-2   -9.955737E-5   -7.252666E-6   7.252666E-6   -9.955737E-5   9.982120E-5   -1.758334E+2   -8.583341E+1   
5.798106E+3   1.967220E+1   1.967220E+1   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   -6.820926E-2   8.893861E-2   -1.000949E-4   -7.695863E-6   7.695863E-6   -1.000949E-4   1.003903E-4   -1.756034E+2   -8.560343E+1   
5.819941E+3   1.965991E+1   1.965991E+1   2.700000E+1   2.700000E+1   9.000000E+1   2.700000E+1   2.700000E+1   -6.826049E-2   8.877416E-2   -1.000195E-4   -7.550455E-6   7.550455E-6   -1.000195E-4   1.003041E-4   -1.756829E+2   -8.568294E+1   
5.842019E+3   1.964910E+1   1.964910E+1   2.900000E+1   2.900000E+1   9.000000E+1   2.900000E+1   2.900000E+1   -6.765978E-2   9.007527E-2   -1.004955E-4   -8.845388E-6   8.845388E-6   -1.004955E-4   1.008840E-4   -1.749699E+2   -8.496992E+1   
5.864113E+3   1.963510E+1   1.963510E+1   3.100000E+1   3.100000E+1   9.000000E+1   3.200000E+1   3.200000E+1   -6.867741E-2   8.892847E-2   -1.003778E-4   -7.342978E-6   7.342978E-6   -1.003778E-4   1.006460E-4   -1.758161E+2   -8.581607E+1   
5.886184E+3   1.962530E+1   1.962530E+1   3.300000E+1   3.300000E+1   9.000000E+1   3.300000E+1   3.300000E+1   -6.741557E-2   8.948713E-2   -9.996148E-5   -8.641506E-6   8.641506E-6   -9.996148E-5   1.003343E-4   -1.750592E+2   -8.505916E+1   
5.908257E+3   1.963781E+1   1.963781E+1   3.500000E+1   3.500000E+1   9.000000E+1   3.500000E+1   3.500000E+1   -6.814910E-2   8.916133E-2   -1.002028E-4   -7.885966E-6   7.885966E-6   -1.002028E-4   1.005126E-4   -1.755001E+2   -8.550009E+1   
5.930372E+3   1.964449E+1   1.964449E+1   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   -6.833472E-2   9.026180E-2   -1.010343E-4   -8.468133E-6   8.468133E-6   -1.010343E-4   1.013885E-4   -1.752090E+2   -8.520898E+1   
5.952253E+3   1.963220E+1   1.963220E+1   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   -6.828257E-2   8.964731E-2   -1.006018E-4   -8.104964E-6   8.104964E-6   -1.006018E-4   1.009278E-4   -1.753939E+2   -8.539393E+1   
5.974189E+3   1.963879E+1   1.963879E+1   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   -6.797026E-2   8.988996E-2   -1.005668E-4   -8.494603E-6   8.494603E-6   -1.005668E-4   1.009249E-4   -1.751718E+2   -8.517184E+1   
5.996079E+3   1.962390E+1   1.962390E+1   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   -6.645070E-2   9.014432E-2   -9.979297E-5   -9.784805E-6   9.784805E-6   -9.979297E-5   1.002715E-4   -1.744000E+2   -8.439999E+1   
6.017954E+3   1.962679E+1   1.962679E+1   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   -6.810953E-2   8.969269E-2   -1.005244E-4   -8.262625E-6   8.262625E-6   -1.005244E-4   1.008634E-4   -1.753011E+2   -8.530112E+1   
6.039805E+3   1.963171E+1   1.963171E+1   4.700000E+1   4.700000E+1   9.000000E+1   4.700000E+1   4.700000E+1   -6.908085E-2   8.946628E-2   -1.009775E-4   -7.396188E-6   7.396188E-6   -1.009775E-4   1.012480E-4   -1.758108E+2   -8.581080E+1   
6.061865E+3   1.962969E+1   1.962969E+1   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   -6.835743E-2   9.092664E-2   -1.014813E-4   -8.885990E-6   8.885990E-6   -1.014813E-4   1.018696E-4   -1.749958E+2   -8.499578E+1   
6.095796E+3   1.962771E+1   1.962771E+1   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   -6.902348E-2   9.110119E-2   -1.020068E-4   -8.507480E-6   8.507480E-6   -1.020068E-4   1.023609E-4   -1.752325E+2   -8.523250E+1   
6.118381E+3   1.962460E+1   1.962460E+1   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   -6.948305E-2   9.335868E-2   -1.037612E-4   -9.643444E-6   9.643444E-6   -1.037612E-4   1.042084E-4   -1.746903E+2   -8.469025E+1   
6.140698E+3   1.962841E+1   1.962841E+1   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   -7.146031E-2   9.342372E-2   -1.050260E-4   -8.223524E-6   8.223524E-6   -1.050260E-4   1.053474E-4   -1.755229E+2   -8.552288E+1   
6.163082E+3   1.962899E+1   1.962899E+1   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   -7.132195E-2   9.499552E-2   -1.059641E-4   -9.353453E-6   9.353453E-6   -1.059641E-4   1.063762E-4   -1.749556E+2   -8.495558E+1   
6.185721E+3   1.961990E+1   1.961990E+1   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   -7.251325E-2   9.589291E-2   -1.072851E-4   -9.059027E-6   9.059027E-6   -1.072851E-4   1.076669E-4   -1.751735E+2   -8.517346E+1   
6.207908E+3   1.960131E+1   1.960131E+1   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   -7.483811E-2   9.745921E-2   -1.097426E-4   -8.363487E-6   8.363487E-6   -1.097426E-4   1.100608E-4   -1.756419E+2   -8.564191E+1   
6.230287E+3   1.961111E+1   1.961111E+1   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   -7.314586E-2   9.900573E-2   -1.097036E-4   -1.062620E-5   1.062620E-5   -1.097036E-4   1.102170E-4   -1.744674E+2   -8.446743E+1   
6.252915E+3   1.962310E+1   1.962310E+1   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   -7.547010E-2   1.001292E-1   -1.118722E-4   -9.641625E-6   9.641625E-6   -1.118722E-4   1.122870E-4   -1.750742E+2   -8.507418E+1   
6.275220E+3   1.961279E+1   1.961279E+1   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   -7.514490E-2   1.014202E-1   -1.125120E-4   -1.072616E-5   1.072616E-5   -1.125120E-4   1.130221E-4   -1.745543E+2   -8.455425E+1   
6.297439E+3   1.962109E+1   1.962109E+1   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   -7.676814E-2   1.023372E-1   -1.141128E-4   -1.012507E-5   1.012507E-5   -1.141128E-4   1.145611E-4   -1.749295E+2   -8.492950E+1   
6.320287E+3   1.961691E+1   1.961691E+1   5.980000E+2   5.980000E+2   9.000000E+1   5.990000E+2   5.990000E+2   -7.682858E-2   1.038181E-1   -1.151146E-4   -1.104853E-5   1.104853E-5   -1.151146E-4   1.156436E-4   -1.745176E+2   -8.451763E+1   
6.342875E+3   1.960281E+1   1.960281E+1   6.480000E+2   6.480000E+2   9.000000E+1   6.480000E+2   6.480000E+2   -7.775171E-2   1.049333E-1   -1.164117E-4   -1.109483E-5   1.109483E-5   -1.164117E-4   1.169392E-4   -1.745558E+2   -8.455576E+1   
6.365516E+3   1.960659E+1   1.960659E+1   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   -7.897182E-2   1.063197E-1   -1.180689E-4   -1.109878E-5   1.109878E-5   -1.180689E-4   1.185895E-4   -1.746298E+2   -8.462983E+1   
6.388921E+3   1.960629E+1   1.960629E+1   7.480000E+2   7.480000E+2   9.000000E+1   7.490000E+2   7.490000E+2   -7.960690E-2   1.073474E-1   -1.191310E-4   -1.130098E-5   1.130098E-5   -1.191310E-4   1.196658E-4   -1.745810E+2   -8.458103E+1   
6.411444E+3   1.959509E+1   1.959509E+1   7.980000E+2   7.980000E+2   9.000000E+1   7.990000E+2   7.990000E+2   -7.877795E-2   1.094462E-1   -1.199854E-4   -1.328622E-5   1.328622E-5   -1.199854E-4   1.207187E-4   -1.736813E+2   -8.368127E+1   
6.433994E+3   1.958599E+1   1.958599E+1   8.480000E+2   8.480000E+2   9.000000E+1   8.480000E+2   8.480000E+2   -8.038276E-2   1.112729E-1   -1.221672E-4   -1.329346E-5   1.329346E-5   -1.221672E-4   1.228883E-4   -1.737899E+2   -8.378987E+1   
6.457352E+3   1.957409E+1   1.957409E+1   8.980000E+2   8.980000E+2   9.000000E+1   8.980000E+2   8.980000E+2   -8.122463E-2   1.121960E-1   -1.232889E-4   -1.327430E-5   1.327430E-5   -1.232889E-4   1.240015E-4   -1.738547E+2   -8.385474E+1   
6.479995E+3   1.956310E+1   1.956310E+1   9.480000E+2   9.480000E+2   9.000000E+1   9.480000E+2   9.480000E+2   -8.238458E-2   1.143184E-1   -1.253883E-4   -1.380393E-5   1.380393E-5   -1.253883E-4   1.261459E-4   -1.737176E+2   -8.371764E+1   
6.502536E+3   1.957672E+1   1.957672E+1   9.980000E+2   9.980000E+2   9.000000E+1   9.990000E+2   9.990000E+2   -8.223947E-2   1.148264E-1   -1.256295E-4   -1.424340E-5   1.424340E-5   -1.256295E-4   1.264344E-4   -1.735316E+2   -8.353164E+1   
6.526078E+3   1.956481E+1   1.956481E+1   1.048000E+3   1.048000E+3   9.000000E+1   1.049000E+3   1.049000E+3   -8.335497E-2   1.162404E-1   -1.272401E-4   -1.434278E-5   1.434278E-5   -1.272401E-4   1.280459E-4   -1.735686E+2   -8.356864E+1   
6.548865E+3   1.956039E+1   1.956039E+1   1.098000E+3   1.098000E+3   9.000000E+1   1.099000E+3   1.099000E+3   -8.475549E-2   1.164343E-1   -1.282322E-4   -1.343368E-5   1.343368E-5   -1.282322E-4   1.289340E-4   -1.740195E+2   -8.401948E+1   
6.571396E+3   1.954949E+1   1.954949E+1   1.148000E+3   1.148000E+3   9.000000E+1   1.149000E+3   1.149000E+3   -8.644469E-2   1.179425E-1   -1.302589E-4   -1.317031E-5   1.317031E-5   -1.302589E-4   1.309230E-4   -1.742265E+2   -8.422652E+1   
6.594456E+3   1.954769E+1   1.954769E+1   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   -8.653120E-2   1.201990E-1   -1.317820E-4   -1.458153E-5   1.458153E-5   -1.317820E-4   1.325862E-4   -1.736860E+2   -8.368597E+1   
6.616991E+3   1.954199E+1   1.954199E+1   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   -8.700612E-2   1.216903E-1   -1.330469E-4   -1.520525E-5   1.520525E-5   -1.330469E-4   1.339129E-4   -1.734802E+2   -8.348024E+1   
6.639578E+3   1.952831E+1   1.952831E+1   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   -8.750895E-2   1.214528E-1   -1.332031E-4   -1.467809E-5   1.467809E-5   -1.332031E-4   1.340093E-4   -1.737118E+2   -8.371176E+1   
6.662607E+3   1.954070E+1   1.954070E+1   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   -8.768443E-2   1.244315E-1   -1.352515E-4   -1.649566E-5   1.649566E-5   -1.352515E-4   1.362537E-4   -1.730464E+2   -8.304638E+1   
6.685177E+3   1.953951E+1   1.953951E+1   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   -8.857752E-2   1.256893E-1   -1.366229E-4   -1.665745E-5   1.665745E-5   -1.366229E-4   1.376346E-4   -1.730486E+2   -8.304865E+1   
6.707687E+3   1.953051E+1   1.953051E+1   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   -8.947396E-2   1.270402E-1   -1.380569E-4   -1.687755E-5   1.687755E-5   -1.380569E-4   1.390847E-4   -1.730301E+2   -8.303014E+1   
6.730483E+3   1.952590E+1   1.952590E+1   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   -9.100734E-2   1.281348E-1   -1.397178E-4   -1.645905E-5   1.645905E-5   -1.397178E-4   1.406839E-4   -1.732814E+2   -8.328140E+1   
6.753028E+3   1.952520E+1   1.952520E+1   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   -9.220049E-2   1.288134E-1   -1.408975E-4   -1.602022E-5   1.602022E-5   -1.408975E-4   1.418053E-4   -1.735133E+2   -8.351326E+1   
6.775559E+3   1.953329E+1   1.953329E+1   1.599000E+3   1.599000E+3   9.000000E+1   1.599000E+3   1.599000E+3   -9.246985E-2   1.311331E-1   -1.425748E-4   -1.733753E-5   1.733753E-5   -1.425748E-4   1.436250E-4   -1.730667E+2   -8.306670E+1   
6.798349E+3   1.953188E+1   1.953188E+1   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   -9.300341E-2   1.315570E-1   -1.431808E-4   -1.722007E-5   1.722007E-5   -1.431808E-4   1.442126E-4   -1.731421E+2   -8.314209E+1   
6.820898E+3   1.952551E+1   1.952551E+1   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   -9.558520E-2   1.334110E-1   -1.459844E-4   -1.652257E-5   1.652257E-5   -1.459844E-4   1.469165E-4   -1.735427E+2   -8.354272E+1   
6.843436E+3   1.954351E+1   1.954351E+1   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   -9.503389E-2   1.346529E-1   -1.464524E-4   -1.774225E-5   1.774225E-5   -1.464524E-4   1.475232E-4   -1.730925E+2   -8.309246E+1   
6.866185E+3   1.954281E+1   1.954281E+1   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   -9.487399E-2   1.359098E-1   -1.471722E-4   -1.868226E-5   1.868226E-5   -1.471722E-4   1.483532E-4   -1.727655E+2   -8.276548E+1   
6.888764E+3   1.953079E+1   1.953079E+1   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   -9.761686E-2   1.373290E-1   -1.497923E-4   -1.758139E-5   1.758139E-5   -1.497923E-4   1.508205E-4   -1.733057E+2   -8.330572E+1   
6.911295E+3   1.952731E+1   1.952731E+1   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   -9.578035E-2   1.381638E-1   -1.492005E-4   -1.948549E-5   1.948549E-5   -1.492005E-4   1.504676E-4   -1.725593E+2   -8.255932E+1   
6.934087E+3   1.953579E+1   1.953579E+1   1.949000E+3   1.949000E+3   9.000000E+1   1.949000E+3   1.949000E+3   -9.766258E-2   1.407001E-1   -1.520160E-4   -1.975146E-5   1.975146E-5   -1.520160E-4   1.532938E-4   -1.725970E+2   -8.259703E+1   
6.956620E+3   1.953430E+1   1.953430E+1   1.999000E+3   1.999000E+3   9.000000E+1   2.000000E+3   2.000000E+3   -9.814883E-2   1.403961E-1   -1.521187E-4   -1.919306E-5   1.919306E-5   -1.521187E-4   1.533247E-4   -1.728089E+2   -8.280890E+1   
6.994566E+3   1.952969E+1   1.952969E+1   2.498000E+3   2.498000E+3   9.000000E+1   2.498000E+3   2.498000E+3   -1.073201E-1   1.551098E-1   -1.673717E-4   -2.202912E-5   2.202912E-5   -1.673717E-4   1.688152E-4   -1.725019E+2   -8.250195E+1   
7.021227E+3   1.953530E+1   1.953530E+1   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   -1.152056E-1   1.688768E-1   -1.812132E-4   -2.519725E-5   2.519725E-5   -1.812132E-4   1.829566E-4   -1.720839E+2   -8.208392E+1   
7.047166E+3   1.952819E+1   1.952819E+1   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -1.253396E-1   1.849111E-1   -1.979214E-4   -2.818460E-5   2.818460E-5   -1.979214E-4   1.999181E-4   -1.718954E+2   -8.189540E+1   
7.073016E+3   1.952831E+1   1.952831E+1   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -1.322743E-1   1.989865E-1   -2.113760E-4   -3.225755E-5   3.225755E-5   -2.113760E-4   2.138232E-4   -1.713232E+2   -8.132318E+1   
7.099677E+3   1.953329E+1   1.953329E+1   4.498000E+3   4.498000E+3   9.000000E+1   4.499000E+3   4.499000E+3   -1.405228E-1   2.133042E-1   -2.258005E-4   -3.551725E-5   3.551725E-5   -2.258005E-4   2.285768E-4   -1.710609E+2   -8.106091E+1   
7.125644E+3   1.949691E+1   1.949691E+1   4.998000E+3   4.998000E+3   9.000000E+1   4.999000E+3   4.999000E+3   -1.480017E-1   2.270169E-1   -2.393553E-4   -3.895054E-5   3.895054E-5   -2.393553E-4   2.425038E-4   -1.707572E+2   -8.075722E+1   
7.151385E+3   1.950460E+1   1.950460E+1   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -1.519379E-1   2.343041E-1   -2.465349E-4   -4.080344E-5   4.080344E-5   -2.465349E-4   2.498887E-4   -1.706023E+2   -8.060230E+1   
7.177835E+3   1.947421E+1   1.947421E+1   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -1.494464E-1   2.368754E-1   -2.466692E-4   -4.432721E-5   4.432721E-5   -2.466692E-4   2.506204E-4   -1.698125E+2   -7.981251E+1   
7.203736E+3   1.949001E+1   1.949001E+1   6.498000E+3   6.498000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -1.397423E-1   2.288932E-1   -2.354709E-4   -4.628620E-5   4.628620E-5   -2.354709E-4   2.399770E-4   -1.688792E+2   -7.887923E+1   
7.229631E+3   1.947000E+1   1.947000E+1   6.998000E+3   6.998000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -1.251221E-1   2.129041E-1   -2.160185E-4   -4.664652E-5   4.664652E-5   -2.160185E-4   2.209975E-4   -1.678148E+2   -7.781478E+1   
7.255332E+3   1.945260E+1   1.945260E+1   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -1.055957E-1   1.942778E-1   -1.918152E-4   -4.891148E-5   4.891148E-5   -1.918152E-4   1.979531E-4   -1.656948E+2   -7.569484E+1   
7.280726E+3   1.946859E+1   1.946859E+1   7.999000E+3   7.999000E+3   9.000000E+1   8.000000E+3   8.000000E+3   -9.077946E-2   1.798336E-1   -1.732478E-4   -5.042682E-5   5.042682E-5   -1.732478E-4   1.804374E-4   -1.637714E+2   -7.377143E+1   
7.307187E+3   1.945721E+1   1.945721E+1   8.498000E+3   8.498000E+3   9.000000E+1   8.499000E+3   8.499000E+3   -8.255059E-2   1.728544E-1   -1.636149E-4   -5.195034E-5   5.195034E-5   -1.636149E-4   1.716644E-4   -1.623845E+2   -7.238452E+1   
7.333555E+3   1.944769E+1   1.944769E+1   8.998000E+3   8.998000E+3   9.000000E+1   8.999000E+3   8.999000E+3   -8.376455E-2   1.778309E-1   -1.676065E-4   -5.430594E-5   5.430594E-5   -1.676065E-4   1.761848E-4   -1.620472E+2   -7.204724E+1   
7.359694E+3   1.945910E+1   1.945910E+1   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -8.882790E-2   1.866802E-1   -1.765004E-4   -5.634638E-5   5.634638E-5   -1.765004E-4   1.852763E-4   -1.622947E+2   -7.229472E+1   
7.384875E+3   1.944521E+1   1.944521E+1   9.999000E+3   9.999000E+3   9.000000E+1   1.000000E+4   1.000000E+4   -9.875900E-2   2.013589E-1   -1.922004E-4   -5.859755E-5   5.859755E-5   -1.922004E-4   2.009344E-4   -1.630447E+2   -7.304472E+1   
@@END Data.
@Time at end of measurement: 12:46:46
@NO Instrument  Changes.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -9499.000      -9998.000      249.500        Coercive Field: Field at which M//H changes sign
Ms  emu                                 3.318E-4       -3.123E-4      3.221E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -9.873E-5      1.515E-4       1.251E-4       Remanent Magnetization: M at H=0        
S                                       0.298          0.485          0.391          Squareness: Mr/Ms                       
S*                                      1.343          1.272          1.307          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
