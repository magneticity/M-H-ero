@Filename: c:\vsm-lv\Will\data\AJA1810b_Pt_CoFeB_Ir8\AJA1810b_Pt_CoFeB_Ir8_OoP_fine.VHD
@Measurement Controlfilename: c:\vsm-lv\Will\Recipes\6_kOe outOfPlane loop (RT).VHC
@Signal Manipulation filename: C:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA1810b_Pt_CoFeB_Ir8
@Date: 18 November 2024    (2024-18-11)
@Time: 18:57:58
@Test ID: 
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 89.9991 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Applied Field to 5999.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Auto Range Signal to 10.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 4
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 10.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 6000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 100.0000 [Oe] Max Stepsize/Sweeprate = 100.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =   10.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To:  0.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =   10.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From:  0.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 10.0000 [Oe] Max Stepsize/Sweeprate = 10.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =   10.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -6000.0000 [Oe] Min Stepsize/Sweeprate = 100.0000 [Oe] Max Stepsize/Sweeprate = 100.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =   10.00 [sec] Up & Down = No
@Section 3 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 5 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.538
@Y Coils Correction Factor: 0.969
@Sample Shape Correction Factor: 0.928
@Coil Angle Alpha: 46.000
@Coil Angle Beta: -43.440
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
14999.000000   1.000000
15248.000000   0.999857
15498.000000   0.999857
15748.000000   0.999857
15999.000000   0.999857
16248.000000   0.999857
16498.000000   0.999857
16748.000000   0.999857
16998.000000   0.999710
17248.000000   0.999710
17498.000000   0.999857
17748.000000   0.999710
17998.000000   0.999857
18248.000000   0.999857
18498.000000   0.999857
18747.000000   0.999710
18997.000000   0.999857
19247.000000   0.999857
19498.000000   0.999857
19748.000000   0.999857
19998.000000   1.000000
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = Yes   Method = Angle Dependent Straight Line
Angular BG Signal array length = 25
Angle = 0.000000, Ofx = 5.511961E-6, Ofy = 7.255357E-5, Ofz = 0.000000E+0,Sx = -6.637759E-8, Sy = 3.436505E-9, Sz = 0.000000E+0
Angle = 15.000000, Ofx = 2.427508E-5, Ofy = 6.341217E-5, Ofz = 0.000000E+0,Sx = -6.122584E-8, Sy = 5.840215E-9, Sz = 0.000000E+0
Angle = 30.000000, Ofx = 3.849872E-5, Ofy = 5.614447E-5, Ofz = 0.000000E+0,Sx = -5.635123E-8, Sy = 5.018955E-9, Sz = 0.000000E+0
Angle = 45.000000, Ofx = 5.162249E-5, Ofy = 4.202634E-5, Ofz = 0.000000E+0,Sx = -5.340771E-8, Sy = 2.320584E-9, Sz = 0.000000E+0
Angle = 60.000000, Ofx = 5.888400E-5, Ofy = 2.821182E-5, Ofz = 0.000000E+0,Sx = -5.406333E-8, Sy = -1.140501E-9, Sz = 0.000000E+0
Angle = 75.000000, Ofx = 6.221306E-5, Ofy = 1.289058E-5, Ofz = 0.000000E+0,Sx = -5.702493E-8, Sy = -3.657483E-9, Sz = 0.000000E+0
Angle = 90.000000, Ofx = 6.528234E-5, Ofy = -3.469610E-6, Ofz = 0.000000E+0,Sx = -6.107239E-8, Sy = -4.959955E-9, Sz = 0.000000E+0
Angle = 105.000000, Ofx = 6.057411E-5, Ofy = -2.091353E-5, Ofz = 0.000000E+0,Sx = -6.580139E-8, Sy = -4.363769E-9, Sz = 0.000000E+0
Angle = 120.000000, Ofx = 5.108214E-5, Ofy = -3.497132E-5, Ofz = 0.000000E+0,Sx = -6.884862E-8, Sy = -3.031072E-9, Sz = 0.000000E+0
Angle = 135.000000, Ofx = 4.040625E-5, Ofy = -4.776267E-5, Ofz = 0.000000E+0,Sx = -7.079075E-8, Sy = -1.151461E-9, Sz = 0.000000E+0
Angle = 150.000000, Ofx = 2.815022E-5, Ofy = -5.275402E-5, Ofz = 0.000000E+0,Sx = -7.120194E-8, Sy = 2.952987E-10, Sz = 0.000000E+0
Angle = 165.000000, Ofx = 1.212763E-5, Ofy = -5.879891E-5, Ofz = 0.000000E+0,Sx = -6.933078E-8, Sy = 2.280793E-9, Sz = 0.000000E+0
Angle = 180.000000, Ofx = -1.503896E-6, Ofy = -5.933596E-5, Ofz = 0.000000E+0,Sx = -6.651357E-8, Sy = 4.300089E-9, Sz = 0.000000E+0
Angle = 195.000000, Ofx = -1.730048E-5, Ofy = -5.754707E-5, Ofz = 0.000000E+0,Sx = -6.233355E-8, Sy = 8.012817E-9, Sz = 0.000000E+0
Angle = 210.000000, Ofx = -3.045760E-5, Ofy = -5.052679E-5, Ofz = 0.000000E+0,Sx = -5.781798E-8, Sy = 6.626921E-9, Sz = 0.000000E+0
Angle = 225.000000, Ofx = -4.215979E-5, Ofy = -4.022672E-5, Ofz = 0.000000E+0,Sx = -5.424357E-8, Sy = 3.244164E-9, Sz = 0.000000E+0
Angle = 240.000000, Ofx = -4.971286E-5, Ofy = -2.831545E-5, Ofz = 0.000000E+0,Sx = -5.470668E-8, Sy = 5.438258E-11, Sz = 0.000000E+0
Angle = 255.000000, Ofx = -5.636146E-5, Ofy = -1.346311E-5, Ofz = 0.000000E+0,Sx = -5.652969E-8, Sy = -2.877288E-9, Sz = 0.000000E+0
Angle = 270.000000, Ofx = -5.608366E-5, Ofy = 3.241239E-6, Ofz = 0.000000E+0,Sx = -6.052403E-8, Sy = -4.749283E-9, Sz = 0.000000E+0
Angle = 285.000000, Ofx = -5.288340E-5, Ofy = 1.695085E-5, Ofz = 0.000000E+0,Sx = -6.466049E-8, Sy = -5.255801E-9, Sz = 0.000000E+0
Angle = 300.000000, Ofx = -4.592161E-5, Ofy = 3.148083E-5, Ofz = 0.000000E+0,Sx = -6.903811E-8, Sy = -4.123988E-9, Sz = 0.000000E+0
Angle = 315.000000, Ofx = -3.562648E-5, Ofy = 4.183753E-5, Ofz = 0.000000E+0,Sx = -7.195187E-8, Sy = -1.570295E-9, Sz = 0.000000E+0
Angle = 330.000000, Ofx = -2.158101E-5, Ofy = 4.883870E-5, Ofz = 0.000000E+0,Sx = -7.205703E-8, Sy = 1.349250E-9, Sz = 0.000000E+0
Angle = 345.000000, Ofx = -8.527411E-6, Ofy = 5.632367E-5, Ofz = 0.000000E+0,Sx = -7.020069E-8, Sy = 3.857333E-9, Sz = 0.000000E+0
Angle = 360.000000, Ofx = 4.810742E-6, Ofy = 5.580095E-5, Ofz = 0.000000E+0,Sx = -6.573828E-8, Sy = 6.096652E-9, Sz = 0.000000E+0
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 15 October 2024  12:22:06
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 4
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 18:57:58
@@Data
New Section: Section 0: 
3.724100E+1   2.064599E+1   2.064599E+1   5.998000E+3   5.998000E+3   8.999910E+1   5.999000E+3   5.999000E+3   4.158982E-2   -3.873698E-2   3.527851E-4   3.157553E-5   -3.156998E-5   3.527856E-4   3.541954E-4   5.114548E+0   9.511365E+1   
6.468800E+1   2.065310E+1   2.065310E+1   5.898000E+3   5.898000E+3   8.999910E+1   5.899000E+3   5.899000E+3   4.778797E-2   -4.280746E-2   3.533301E-4   2.963669E-5   -2.963114E-5   3.533306E-4   3.545709E-4   4.794642E+0   9.479374E+1   
9.214800E+1   2.066259E+1   2.066259E+1   5.798000E+3   5.798000E+3   8.999910E+1   5.799000E+3   5.799000E+3   5.346262E-2   -4.950044E-2   3.551462E-4   2.990584E-5   -2.990026E-5   3.551467E-4   3.564031E-4   4.813357E+0   9.481246E+1   
1.193660E+2   2.064980E+1   2.064980E+1   5.698000E+3   5.698000E+3   8.999910E+1   5.699000E+3   5.699000E+3   5.707753E-2   -5.340366E-2   3.538636E-4   2.964381E-5   -2.963826E-5   3.538641E-4   3.551031E-4   4.788593E+0   9.478769E+1   
1.468230E+2   2.063339E+1   2.063339E+1   5.599000E+3   5.599000E+3   8.999910E+1   5.599000E+3   5.599000E+3   6.064055E-2   -5.969315E-2   3.540209E-4   3.109605E-5   -3.109049E-5   3.540214E-4   3.553840E-4   5.019791E+0   9.501889E+1   
1.749710E+2   2.063061E+1   2.063061E+1   5.498000E+3   5.498000E+3   8.999910E+1   5.499000E+3   5.499000E+3   6.743283E-2   -6.431476E-2   3.553030E-4   2.913209E-5   -2.912651E-5   3.553035E-4   3.564953E-4   4.687325E+0   9.468642E+1   
2.021710E+2   2.062670E+1   2.062670E+1   5.398000E+3   5.398000E+3   8.999910E+1   5.399000E+3   5.399000E+3   7.119075E-2   -6.873726E-2   3.544368E-4   2.913592E-5   -2.913036E-5   3.544373E-4   3.556323E-4   4.699344E+0   9.469844E+1   
2.296190E+2   2.062689E+1   2.062689E+1   5.298000E+3   5.298000E+3   8.999910E+1   5.299000E+3   5.299000E+3   7.695671E-2   -7.488237E-2   3.559753E-4   2.895634E-5   -2.895075E-5   3.559757E-4   3.571510E-4   4.650412E+0   9.464951E+1   
2.571100E+2   2.061450E+1   2.061450E+1   5.198000E+3   5.198000E+3   8.999910E+1   5.199000E+3   5.199000E+3   8.189706E-2   -7.876640E-2   3.555655E-4   2.776011E-5   -2.775452E-5   3.555659E-4   3.566475E-4   4.464205E+0   9.446330E+1   
2.842960E+2   2.060479E+1   2.060479E+1   5.098000E+3   5.098000E+3   8.999910E+1   5.099000E+3   5.099000E+3   8.680674E-2   -8.360337E-2   3.557241E-4   2.725535E-5   -2.724976E-5   3.557245E-4   3.567667E-4   4.381405E+0   9.438051E+1   
3.115040E+2   2.059899E+1   2.059899E+1   4.998000E+3   4.998000E+3   8.999910E+1   4.999000E+3   4.999000E+3   9.286347E-2   -8.986771E-2   3.575303E-4   2.695765E-5   -2.695203E-5   3.575307E-4   3.585452E-4   4.311920E+0   9.431102E+1   
3.387200E+2   2.059271E+1   2.059271E+1   4.898000E+3   4.898000E+3   8.999910E+1   4.899000E+3   4.899000E+3   9.851525E-2   -9.524696E-2   3.585193E-4   2.631878E-5   -2.631314E-5   3.585198E-4   3.594841E-4   4.198531E+0   9.419763E+1   
3.675510E+2   2.058090E+1   2.058090E+1   4.798000E+3   4.798000E+3   8.999910E+1   4.799000E+3   4.799000E+3   1.027700E-1   -9.893350E-2   3.575299E-4   2.545991E-5   -2.545429E-5   3.575303E-4   3.584353E-4   4.073189E+0   9.407229E+1   
3.947240E+2   2.057980E+1   2.057980E+1   4.698000E+3   4.698000E+3   8.999910E+1   4.699000E+3   4.699000E+3   1.073279E-1   -1.054600E-1   3.584977E-4   2.638776E-5   -2.638213E-5   3.584981E-4   3.594676E-4   4.209749E+0   9.420885E+1   
4.221200E+2   2.058099E+1   2.058099E+1   4.598000E+3   4.598000E+3   8.999910E+1   4.599000E+3   4.599000E+3   1.131939E-1   -1.107393E-1   3.595680E-4   2.552971E-5   -2.552406E-5   3.595684E-4   3.604732E-4   4.061247E+0   9.406035E+1   
4.493500E+2   2.057189E+1   2.057189E+1   4.498000E+3   4.498000E+3   8.999910E+1   4.499000E+3   4.499000E+3   1.167586E-1   -1.142183E-1   3.579898E-4   2.500425E-5   -2.499862E-5   3.579902E-4   3.588620E-4   3.995407E+0   9.399451E+1   
4.768220E+2   2.056130E+1   2.056130E+1   4.399000E+3   4.399000E+3   8.999910E+1   4.399000E+3   4.399000E+3   1.219827E-1   -1.200801E-1   3.589915E-4   2.500188E-5   -2.499624E-5   3.589919E-4   3.598611E-4   3.983918E+0   9.398302E+1   
5.042970E+2   2.054449E+1   2.054449E+1   4.299000E+3   4.299000E+3   8.999910E+1   4.299000E+3   4.299000E+3   1.273987E-1   -1.272186E-1   3.609102E-4   2.576400E-5   -2.575833E-5   3.609106E-4   3.618287E-4   4.083200E+0   9.408230E+1   
5.314920E+2   2.054821E+1   2.054821E+1   4.199000E+3   4.199000E+3   8.999910E+1   4.199000E+3   4.199000E+3   1.316686E-1   -1.317641E-1   3.604617E-4   2.549868E-5   -2.549302E-5   3.604621E-4   3.613625E-4   4.046303E+0   9.404540E+1   
5.592440E+2   2.053619E+1   2.053619E+1   4.099000E+3   4.099000E+3   8.999910E+1   4.100000E+3   4.100000E+3   1.390687E-1   -1.362399E-1   3.621204E-4   2.301491E-5   -2.300922E-5   3.621208E-4   3.628510E-4   3.636596E+0   9.363570E+1   
5.869040E+2   2.053439E+1   2.053439E+1   3.999000E+3   3.999000E+3   8.999910E+1   4.000000E+3   4.000000E+3   1.436066E-1   -1.421863E-1   3.627165E-4   2.354871E-5   -2.354302E-5   3.627168E-4   3.634801E-4   3.714612E+0   9.371371E+1   
6.145040E+2   2.053860E+1   2.053860E+1   3.899000E+3   3.899000E+3   8.999910E+1   3.900000E+3   3.900000E+3   1.483312E-1   -1.460338E-1   3.621401E-4   2.247656E-5   -2.247087E-5   3.621405E-4   3.628370E-4   3.551560E+0   9.355066E+1   
6.421230E+2   2.052249E+1   2.052249E+1   3.799000E+3   3.799000E+3   8.999910E+1   3.800000E+3   3.800000E+3   1.528101E-1   -1.515147E-1   3.624092E-4   2.272393E-5   -2.271824E-5   3.624095E-4   3.631209E-4   3.587886E+0   9.358699E+1   
6.700350E+2   2.054141E+1   2.054141E+1   3.699000E+3   3.699000E+3   8.999910E+1   3.700000E+3   3.700000E+3   1.569338E-1   -1.584513E-1   3.633406E-4   2.424183E-5   -2.423612E-5   3.633409E-4   3.641484E-4   3.817078E+0   9.381618E+1   
6.977100E+2   2.054290E+1   2.054290E+1   3.599000E+3   3.599000E+3   8.999910E+1   3.600000E+3   3.600000E+3   1.608514E-1   -1.606354E-1   3.611978E-4   2.256047E-5   -2.255479E-5   3.611981E-4   3.619016E-4   3.574060E+0   9.357316E+1   
7.257800E+2   2.053729E+1   2.053729E+1   3.499000E+3   3.499000E+3   8.999910E+1   3.499000E+3   3.499000E+3   1.678682E-1   -1.662728E-1   3.631963E-4   2.114999E-5   -2.114428E-5   3.631966E-4   3.638116E-4   3.332738E+0   9.333184E+1   
7.539230E+2   2.054611E+1   2.054611E+1   3.398000E+3   3.398000E+3   8.999910E+1   3.399000E+3   3.399000E+3   1.727137E-1   -1.719101E-1   3.638066E-4   2.125268E-5   -2.124697E-5   3.638069E-4   3.644268E-4   3.343278E+0   9.334238E+1   
7.811100E+2   2.054119E+1   2.054119E+1   3.299000E+3   3.299000E+3   8.999910E+1   3.299000E+3   3.299000E+3   1.782714E-1   -1.783195E-1   3.653694E-4   2.140366E-5   -2.139792E-5   3.653697E-4   3.659958E-4   3.352605E+0   9.335171E+1   
8.083130E+2   2.054180E+1   2.054180E+1   3.199000E+3   3.199000E+3   8.999910E+1   3.199000E+3   3.199000E+3   1.823118E-1   -1.823477E-1   3.644480E-4   2.093398E-5   -2.092825E-5   3.644483E-4   3.650487E-4   3.287471E+0   9.328657E+1   
8.357930E+2   2.053439E+1   2.053439E+1   3.099000E+3   3.099000E+3   8.999910E+1   3.099000E+3   3.099000E+3   1.878996E-1   -1.872963E-1   3.651282E-4   2.003659E-5   -2.003085E-5   3.651285E-4   3.656776E-4   3.140983E+0   9.314008E+1   
8.634510E+2   2.053829E+1   2.053829E+1   2.999000E+3   2.999000E+3   8.999910E+1   2.999000E+3   2.999000E+3   1.917723E-1   -1.938935E-1   3.656824E-4   2.149019E-5   -2.148444E-5   3.656827E-4   3.663133E-4   3.363253E+0   9.336235E+1   
8.915190E+2   2.053710E+1   2.053710E+1   2.899000E+3   2.899000E+3   8.999910E+1   2.899000E+3   2.899000E+3   1.963046E-1   -1.973004E-1   3.647055E-4   2.024180E-5   -2.023607E-5   3.647058E-4   3.652668E-4   3.176758E+0   9.317586E+1   
9.196690E+2   2.054119E+1   2.054119E+1   2.799000E+3   2.799000E+3   8.999910E+1   2.799000E+3   2.799000E+3   2.021571E-1   -2.022773E-1   3.655798E-4   1.918053E-5   -1.917479E-5   3.655801E-4   3.660827E-4   3.003330E+0   9.300243E+1   
9.477690E+2   2.054400E+1   2.054400E+1   2.698000E+3   2.698000E+3   8.999910E+1   2.699000E+3   2.699000E+3   2.059717E-1   -2.076390E-1   3.653317E-4   1.980551E-5   -1.979977E-5   3.653320E-4   3.658682E-4   3.103104E+0   9.310220E+1   
9.759060E+2   2.052911E+1   2.052911E+1   2.598000E+3   2.598000E+3   8.999910E+1   2.599000E+3   2.599000E+3   2.101867E-1   -2.116171E-1   3.644960E-4   1.917933E-5   -1.917361E-5   3.644963E-4   3.650003E-4   3.012055E+0   9.301116E+1   
1.005010E+3   2.052700E+1   2.052700E+1   2.498000E+3   2.498000E+3   8.999910E+1   2.499000E+3   2.499000E+3   2.163616E-1   -2.184240E-1   3.667163E-4   1.918105E-5   -1.917529E-5   3.667166E-4   3.672176E-4   2.994121E+0   9.299322E+1   
1.032659E+3   2.051800E+1   2.051800E+1   2.398000E+3   2.398000E+3   8.999910E+1   2.399000E+3   2.399000E+3   2.215529E-1   -2.224917E-1   3.665875E-4   1.793968E-5   -1.793392E-5   3.665878E-4   3.670262E-4   2.801647E+0   9.280075E+1   
1.060753E+3   2.051339E+1   2.051339E+1   2.299000E+3   2.299000E+3   8.999910E+1   2.299000E+3   2.299000E+3   2.255472E-1   -2.269787E-1   3.659189E-4   1.782468E-5   -1.781893E-5   3.659192E-4   3.663528E-4   2.788793E+0   9.278789E+1   
1.088900E+3   2.050680E+1   2.050680E+1   2.199000E+3   2.199000E+3   8.999910E+1   2.199000E+3   2.199000E+3   2.305388E-1   -2.338732E-1   3.674036E-4   1.871006E-5   -1.870429E-5   3.674039E-4   3.678797E-4   2.915274E+0   9.291437E+1   
1.117011E+3   2.052239E+1   2.052239E+1   2.099000E+3   2.099000E+3   8.999910E+1   2.100000E+3   2.100000E+3   2.345066E-1   -2.380124E-1   3.665635E-4   1.837386E-5   -1.836810E-5   3.665638E-4   3.670237E-4   2.869528E+0   9.286863E+1   
1.145573E+3   2.052041E+1   2.052041E+1   1.999000E+3   1.999000E+3   8.999910E+1   2.000000E+3   2.000000E+3   2.392258E-1   -2.396928E-1   3.646444E-4   1.578138E-5   -1.577566E-5   3.646447E-4   3.649858E-4   2.478148E+0   9.247725E+1   
1.184546E+3   2.051211E+1   2.051211E+1   1.949000E+3   1.949000E+3   8.999910E+1   1.950000E+3   1.950000E+3   2.414443E-1   -2.433059E-1   3.653042E-4   1.653341E-5   -1.652767E-5   3.653044E-4   3.656781E-4   2.591398E+0   9.259050E+1   
1.212205E+3   2.051269E+1   2.051269E+1   1.899000E+3   1.899000E+3   8.999910E+1   1.899000E+3   1.899000E+3   2.439921E-1   -2.472716E-1   3.663406E-4   1.729960E-5   -1.729384E-5   3.663408E-4   3.667488E-4   2.703654E+0   9.270275E+1   
1.239404E+3   2.050921E+1   2.050921E+1   1.849000E+3   1.849000E+3   8.999910E+1   1.850000E+3   1.850000E+3   2.474438E-1   -2.498298E-1   3.672326E-4   1.645793E-5   -1.645216E-5   3.672329E-4   3.676012E-4   2.566055E+0   9.256516E+1   
1.266797E+3   2.050521E+1   2.050521E+1   1.799000E+3   1.799000E+3   8.999910E+1   1.800000E+3   1.800000E+3   2.487565E-1   -2.541221E-1   3.677075E-4   1.831682E-5   -1.831104E-5   3.677077E-4   3.681634E-4   2.851749E+0   9.285085E+1   
1.294152E+3   2.049911E+1   2.049911E+1   1.749000E+3   1.749000E+3   8.999910E+1   1.749000E+3   1.749000E+3   2.504799E-1   -2.549824E-1   3.662747E-4   1.747171E-5   -1.746596E-5   3.662749E-4   3.666911E-4   2.731003E+0   9.273010E+1   
1.321557E+3   2.048501E+1   2.048501E+1   1.699000E+3   1.699000E+3   8.999910E+1   1.700000E+3   1.700000E+3   2.532481E-1   -2.572283E-1   3.665175E-4   1.688524E-5   -1.687948E-5   3.665178E-4   3.669063E-4   2.637717E+0   9.263682E+1   
1.348953E+3   2.047561E+1   2.047561E+1   1.649000E+3   1.649000E+3   8.999910E+1   1.650000E+3   1.650000E+3   2.550927E-1   -2.588115E-1   3.656734E-4   1.646929E-5   -1.646355E-5   3.656736E-4   3.660441E-4   2.578760E+0   9.257786E+1   
1.376154E+3   2.047799E+1   2.047799E+1   1.599000E+3   1.599000E+3   8.999910E+1   1.600000E+3   1.600000E+3   2.586155E-1   -2.626599E-1   3.673491E-4   1.648068E-5   -1.647491E-5   3.673494E-4   3.677186E-4   2.568784E+0   9.256788E+1   
1.403878E+3   2.047051E+1   2.047051E+1   1.549000E+3   1.549000E+3   8.999910E+1   1.550000E+3   1.550000E+3   2.608560E-1   -2.654503E-1   3.675152E-4   1.663881E-5   -1.663304E-5   3.675155E-4   3.678916E-4   2.592228E+0   9.259133E+1   
1.431530E+3   2.048400E+1   2.048400E+1   1.499000E+3   1.499000E+3   8.999910E+1   1.500000E+3   1.500000E+3   2.644608E-1   -2.662339E-1   3.673518E-4   1.443782E-5   -1.443205E-5   3.673520E-4   3.676354E-4   2.250705E+0   9.224981E+1   
1.458953E+3   2.047350E+1   2.047350E+1   1.449000E+3   1.449000E+3   8.999910E+1   1.449000E+3   1.449000E+3   2.641410E-1   -2.701712E-1   3.664566E-4   1.717606E-5   -1.717030E-5   3.664568E-4   3.668589E-4   2.683527E+0   9.268263E+1   
1.486380E+3   2.046429E+1   2.046429E+1   1.399000E+3   1.399000E+3   8.999910E+1   1.399000E+3   1.399000E+3   2.672413E-1   -2.713025E-1   3.661713E-4   1.557009E-5   -1.556434E-5   3.661716E-4   3.665022E-4   2.434827E+0   9.243393E+1   
1.513726E+3   2.048919E+1   2.048919E+1   1.349000E+3   1.349000E+3   8.999910E+1   1.349000E+3   1.349000E+3   2.699409E-1   -2.747948E-1   3.670775E-4   1.590286E-5   -1.589710E-5   3.670778E-4   3.674218E-4   2.480668E+0   9.247977E+1   
1.541075E+3   2.047900E+1   2.047900E+1   1.299000E+3   1.299000E+3   8.999910E+1   1.299000E+3   1.299000E+3   2.718395E-1   -2.778638E-1   3.671875E-4   1.649438E-5   -1.648861E-5   3.671878E-4   3.675578E-4   2.572046E+0   9.257115E+1   
1.568411E+3   2.048550E+1   2.048550E+1   1.248000E+3   1.248000E+3   8.999910E+1   1.249000E+3   1.249000E+3   2.736912E-1   -2.770507E-1   3.648675E-4   1.438824E-5   -1.438250E-5   3.648677E-4   3.651511E-4   2.258240E+0   9.225734E+1   
1.595723E+3   2.049160E+1   2.049160E+1   1.199000E+3   1.199000E+3   8.999910E+1   1.199000E+3   1.199000E+3   2.743679E-1   -2.808600E-1   3.646193E-4   1.634917E-5   -1.634344E-5   3.646195E-4   3.649856E-4   2.567367E+0   9.256647E+1   
1.622872E+3   2.049151E+1   2.049151E+1   1.148000E+3   1.148000E+3   8.999910E+1   1.149000E+3   1.149000E+3   2.804302E-1   -2.862767E-1   3.689591E-4   1.569951E-5   -1.569371E-5   3.689593E-4   3.692930E-4   2.436512E+0   9.243561E+1   
1.650259E+3   2.048431E+1   2.048431E+1   1.098000E+3   1.098000E+3   8.999910E+1   1.099000E+3   1.099000E+3   2.820113E-1   -2.866308E-1   3.671796E-4   1.460223E-5   -1.459646E-5   3.671798E-4   3.674698E-4   2.277375E+0   9.227647E+1   
1.677615E+3   2.048431E+1   2.048431E+1   1.048000E+3   1.048000E+3   8.999910E+1   1.049000E+3   1.049000E+3   2.814975E-1   -2.881236E-1   3.647055E-4   1.576097E-5   -1.575524E-5   3.647058E-4   3.650459E-4   2.474532E+0   9.247363E+1   
1.704762E+3   2.046581E+1   2.046581E+1   9.980000E+2   9.980000E+2   8.999910E+1   9.990000E+2   9.990000E+2   2.863642E-1   -2.915926E-1   3.670437E-4   1.457201E-5   -1.456624E-5   3.670440E-4   3.673329E-4   2.273506E+0   9.227261E+1   
1.731715E+3   2.047161E+1   2.047161E+1   9.480000E+2   9.480000E+2   8.999910E+1   9.490000E+2   9.490000E+2   2.870590E-1   -2.922939E-1   3.648871E-4   1.433456E-5   -1.432883E-5   3.648874E-4   3.651686E-4   2.249704E+0   9.224880E+1   
1.758633E+3   2.048480E+1   2.048480E+1   8.980000E+2   8.980000E+2   8.999910E+1   8.990000E+2   8.990000E+2   2.660472E-1   -2.685228E-1   3.331206E-4   1.196472E-5   -1.195949E-5   3.331208E-4   3.333354E-4   2.057013E+0   9.205611E+1   
1.785580E+3   2.047790E+1   2.047790E+1   8.480000E+2   8.480000E+2   8.999910E+1   8.490000E+2   8.490000E+2   1.986102E-1   -1.930980E-1   2.384497E-4   5.517014E-6   -5.513268E-6   2.384498E-4   2.385135E-4   1.325417E+0   9.132452E+1   
1.812516E+3   2.047531E+1   2.047531E+1   7.980000E+2   7.980000E+2   8.999910E+1   7.990000E+2   7.990000E+2   1.745454E-1   -1.687059E-1   2.042617E-4   4.831151E-6   -4.827943E-6   2.042618E-4   2.043188E-4   1.354894E+0   9.135399E+1   
1.839468E+3   2.046621E+1   2.046621E+1   7.480000E+2   7.480000E+2   8.999910E+1   7.490000E+2   7.490000E+2   1.574106E-1   -1.539712E-1   1.806665E-4   6.123207E-6   -6.120369E-6   1.806666E-4   1.807703E-4   1.941144E+0   9.194024E+1   
1.866367E+3   2.045471E+1   2.045471E+1   6.980000E+2   6.980000E+2   8.999910E+1   6.990000E+2   6.990000E+2   1.452760E-1   -1.355058E-1   1.581036E-4   1.318217E-6   -1.315733E-6   1.581036E-4   1.581090E-4   4.777028E-1   9.047680E+1   
1.893326E+3   2.044369E+1   2.044369E+1   6.480000E+2   6.480000E+2   8.999910E+1   6.490000E+2   6.490000E+2   1.328388E-1   -1.247624E-1   1.401102E-4   2.154117E-6   -2.151916E-6   1.401102E-4   1.401267E-4   8.808217E-1   9.087992E+1   
1.920271E+3   2.045580E+1   2.045580E+1   5.990000E+2   5.990000E+2   8.999910E+1   5.990000E+2   5.990000E+2   1.230906E-1   -1.159262E-1   1.250900E-4   2.463355E-6   -2.461390E-6   1.250901E-4   1.251143E-4   1.128160E+0   9.112726E+1   
1.947210E+3   2.044811E+1   2.044811E+1   5.480000E+2   5.480000E+2   8.999910E+1   5.490000E+2   5.490000E+2   1.136446E-1   -1.069860E-1   1.102073E-4   2.489532E-6   -2.487801E-6   1.102074E-4   1.102355E-4   1.294065E+0   9.129316E+1   
1.974196E+3   2.046011E+1   2.046011E+1   4.990000E+2   4.990000E+2   8.999910E+1   5.000000E+2   5.000000E+2   1.022415E-1   -9.493099E-2   9.215482E-5   1.689626E-6   -1.688178E-6   9.215484E-5   9.217031E-5   1.050380E+0   9.104948E+1   
2.001251E+3   2.044781E+1   2.044781E+1   4.490000E+2   4.490000E+2   8.999910E+1   4.500000E+2   4.500000E+2   9.591617E-2   -8.921759E-2   8.134894E-5   1.817400E-6   -1.816123E-6   8.134897E-5   8.136924E-5   1.279821E+0   9.127892E+1   
2.028250E+3   2.044860E+1   2.044860E+1   3.990000E+2   3.990000E+2   8.999910E+1   4.000000E+2   4.000000E+2   8.768634E-2   -7.826170E-2   6.603247E-5   -4.187980E-7   4.198352E-7   6.603246E-5   6.603380E-5   -3.633824E-1   8.963572E+1   
2.055251E+3   2.043301E+1   2.043301E+1   3.490000E+2   3.490000E+2   8.999910E+1   3.500000E+2   3.500000E+2   8.357380E-2   -6.152184E-2   4.989007E-5   -9.582805E-6   9.583589E-6   4.988992E-5   5.080206E-5   -1.087286E+1   7.912624E+1   
2.082251E+3   2.043490E+1   2.043490E+1   2.990000E+2   2.990000E+2   8.999910E+1   3.000000E+2   3.000000E+2   7.041109E-2   -6.121711E-2   3.786269E-5   -9.016575E-7   9.022522E-7   3.786267E-5   3.787342E-5   -1.364177E+0   8.863492E+1   
2.109248E+3   2.043090E+1   2.043090E+1   2.490000E+2   2.490000E+2   8.999910E+1   2.500000E+2   2.500000E+2   6.404930E-2   -5.197710E-2   2.485332E-5   -3.228751E-6   3.229141E-6   2.485327E-5   2.506217E-5   -7.401969E+0   8.259713E+1   
2.136290E+3   2.042501E+1   2.042501E+1   1.990000E+2   1.990000E+2   8.999910E+1   2.000000E+2   2.000000E+2   5.621975E-2   -4.806410E-2   1.415594E-5   -7.898895E-7   7.901119E-7   1.415593E-5   1.417796E-5   -3.193743E+0   8.680536E+1   
2.163269E+3   2.042199E+1   2.042199E+1   1.490000E+2   1.490000E+2   8.999910E+1   1.500000E+2   1.500000E+2   5.229095E-2   -4.499973E-2   6.586521E-6   -4.638555E-7   4.639589E-7   6.586513E-6   6.602834E-6   -4.028402E+0   8.597070E+1   
2.190670E+3   2.041070E+1   2.041070E+1   9.900000E+1   9.900000E+1   8.999910E+1   1.000000E+2   1.000000E+2   4.479888E-2   -3.941518E-2   -4.918479E-6   5.650070E-7   -5.650842E-7   -4.918470E-6   4.950825E-6   1.734469E+2   2.634460E+2   
2.217459E+3   2.042669E+1   2.042669E+1   4.900000E+1   4.900000E+1   8.999910E+1   5.000000E+1   5.000000E+1   3.787946E-2   -3.306122E-2   -1.651669E-5   6.549763E-7   -6.552357E-7   -1.651668E-5   1.652967E-5   1.777291E+2   2.677282E+2   
2.243972E+3   2.043920E+1   2.043920E+1   0.000000E+0   0.000000E+0   8.999910E+1   0.000000E+0   0.000000E+0   2.941643E-2   -2.188786E-2   -3.212319E-5   -1.572177E-6   1.571672E-6   -3.212321E-5   3.216164E-5   -1.771981E+2   -8.719896E+1   
2.282220E+3   2.042611E+1   2.042611E+1   -9.000000E+0   -9.000000E+0   8.999910E+1   -8.000000E+0   -8.000000E+0   2.975892E-2   -2.678532E-2   -2.935694E-5   1.594511E-6   -1.594972E-6   -2.935692E-5   2.940021E-5   1.768911E+2   2.668902E+2   
2.308877E+3   2.043011E+1   2.043011E+1   -1.900000E+1   -1.900000E+1   8.999910E+1   -1.800000E+1   -1.800000E+1   2.757147E-2   -2.658298E-2   -3.155271E-5   2.922126E-6   -2.922622E-6   -3.155266E-5   3.168773E-5   1.747089E+2   2.647080E+2   
2.335602E+3   2.043221E+1   2.043221E+1   -2.900000E+1   -2.900000E+1   8.999910E+1   -2.800000E+1   -2.800000E+1   2.662690E-2   -2.375384E-2   -3.454207E-5   1.538993E-6   -1.539535E-6   -3.454204E-5   3.457633E-5   1.774489E+2   2.674480E+2   
2.362280E+3   2.043649E+1   2.043649E+1   -3.900000E+1   -3.900000E+1   8.999910E+1   -3.800000E+1   -3.800000E+1   2.547878E-2   -2.383367E-2   -3.586977E-5   2.343080E-6   -2.343644E-6   -3.586973E-5   3.594622E-5   1.762626E+2   2.662617E+2   
2.388933E+3   2.045300E+1   2.045300E+1   -4.900000E+1   -4.900000E+1   8.999910E+1   -4.800000E+1   -4.800000E+1   2.418502E-2   -2.463230E-2   -3.685053E-5   3.753843E-6   -3.754422E-6   -3.685047E-5   3.704123E-5   1.741835E+2   2.641826E+2   
2.415625E+3   2.044991E+1   2.044991E+1   -5.900000E+1   -5.900000E+1   8.999910E+1   -5.800000E+1   -5.800000E+1   2.217977E-2   -2.120471E-2   -4.091763E-5   2.686640E-6   -2.687283E-6   -4.091758E-5   4.100573E-5   1.762434E+2   2.662425E+2   
2.442267E+3   2.044259E+1   2.044259E+1   -6.900000E+1   -6.900000E+1   8.999910E+1   -6.800000E+1   -6.800000E+1   1.952368E-2   -1.780853E-2   -4.539972E-5   2.093626E-6   -2.094340E-6   -4.539969E-5   4.544797E-5   1.773597E+2   2.673588E+2   
2.468943E+3   2.043990E+1   2.043990E+1   -7.900000E+1   -7.900000E+1   8.999910E+1   -7.800000E+1   -7.800000E+1   1.939784E-2   -1.692399E-2   -4.664101E-5   1.509364E-6   -1.510096E-6   -4.664099E-5   4.666543E-5   1.781465E+2   2.681456E+2   
2.495589E+3   2.043710E+1   2.043710E+1   -8.900000E+1   -8.900000E+1   8.999910E+1   -8.800000E+1   -8.800000E+1   1.789415E-2   -1.648095E-2   -4.852914E-5   2.192725E-6   -2.193487E-6   -4.852910E-5   4.857865E-5   1.774129E+2   2.674120E+2   
2.522253E+3   2.043179E+1   2.043179E+1   -9.900000E+1   -9.900000E+1   8.999910E+1   -9.800000E+1   -9.800000E+1   1.653305E-2   -1.649284E-2   -5.004098E-5   3.096967E-6   -3.097753E-6   -5.004093E-5   5.013672E-5   1.764586E+2   2.664577E+2   
2.549037E+3   2.043310E+1   2.043310E+1   -1.090000E+2   -1.090000E+2   8.999910E+1   -1.080000E+2   -1.080000E+2   1.418900E-2   -1.272917E-2   -5.454188E-5   2.028755E-6   -2.029612E-6   -5.454185E-5   5.457960E-5   1.778698E+2   2.678689E+2   
2.575882E+3   2.042849E+1   2.042849E+1   -1.190000E+2   -1.190000E+2   8.999910E+1   -1.180000E+2   -1.180000E+2   1.424293E-2   -1.177089E-2   -5.570875E-5   1.267758E-6   -1.268633E-6   -5.570873E-5   5.572317E-5   1.786964E+2   2.686955E+2   
2.602679E+3   2.042391E+1   2.042391E+1   -1.290000E+2   -1.290000E+2   8.999910E+1   -1.280000E+2   -1.280000E+2   1.208595E-2   -1.210514E-2   -5.755261E-5   2.951565E-6   -2.952469E-6   -5.755256E-5   5.762824E-5   1.770642E+2   2.670633E+2   
2.629482E+3   2.040859E+1   2.040859E+1   -1.390000E+2   -1.390000E+2   8.999910E+1   -1.380000E+2   -1.380000E+2   1.088238E-2   -1.124041E-2   -5.950099E-5   3.129875E-6   -3.130810E-6   -5.950094E-5   5.958325E-5   1.769889E+2   2.669880E+2   
2.656243E+3   2.040319E+1   2.040319E+1   -1.490000E+2   -1.490000E+2   8.999910E+1   -1.480000E+2   -1.480000E+2   1.002160E-2   -1.135070E-2   -6.061808E-5   3.755785E-6   -3.756737E-6   -6.061803E-5   6.073432E-5   1.764546E+2   2.664537E+2   
2.683087E+3   2.040460E+1   2.040460E+1   -1.590000E+2   -1.590000E+2   8.999910E+1   -1.580000E+2   -1.580000E+2   7.781444E-3   -6.911827E-3   -6.546687E-5   2.140542E-6   -2.141570E-6   -6.546684E-5   6.550186E-5   1.781273E+2   2.681264E+2   
2.709988E+3   2.040621E+1   2.040621E+1   -1.690000E+2   -1.690000E+2   8.999910E+1   -1.680000E+2   -1.680000E+2   7.603802E-3   -6.922489E-3   -6.618957E-5   2.221840E-6   -2.222880E-6   -6.618954E-5   6.622685E-5   1.780774E+2   2.680765E+2   
2.736801E+3   2.039880E+1   2.039880E+1   -1.790000E+2   -1.790000E+2   8.999910E+1   -1.780000E+2   -1.780000E+2   5.855737E-3   -7.777178E-3   -6.743891E-5   3.987616E-6   -3.988675E-6   -6.743885E-5   6.755670E-5   1.766161E+2   2.666152E+2   
2.763611E+3   2.039520E+1   2.039520E+1   -1.890000E+2   -1.890000E+2   8.999910E+1   -1.880000E+2   -1.880000E+2   5.015676E-3   -5.124148E-3   -7.024969E-5   2.655744E-6   -2.656848E-6   -7.024965E-5   7.029987E-5   1.778350E+2   2.678341E+2   
2.790458E+3   2.038760E+1   2.038760E+1   -1.990000E+2   -1.990000E+2   8.999910E+1   -1.980000E+2   -1.980000E+2   3.157917E-3   -2.411094E-3   -7.377682E-5   1.988603E-6   -1.989761E-6   -7.377679E-5   7.380362E-5   1.784560E+2   2.684551E+2   
2.817304E+3   2.039861E+1   2.039861E+1   -2.090000E+2   -2.090000E+2   8.999910E+1   -2.080000E+2   -2.080000E+2   2.684412E-3   -4.732610E-3   -7.326908E-5   3.900594E-6   -3.901745E-6   -7.326902E-5   7.337283E-5   1.769526E+2   2.669517E+2   
2.844144E+3   2.038311E+1   2.038311E+1   -2.190000E+2   -2.190000E+2   8.999910E+1   -2.180000E+2   -2.180000E+2   8.976483E-4   -1.022877E-3   -7.736469E-5   2.483193E-6   -2.484408E-6   -7.736465E-5   7.740453E-5   1.781616E+2   2.681607E+2   
2.870939E+3   2.039700E+1   2.039700E+1   -2.290000E+2   -2.290000E+2   8.999910E+1   -2.280000E+2   -2.280000E+2   -1.112461E-3   -1.916874E-3   -7.876465E-5   4.458641E-6   -4.459878E-6   -7.876458E-5   7.889074E-5   1.767601E+2   2.667592E+2   
2.897783E+3   2.039211E+1   2.039211E+1   -2.390000E+2   -2.390000E+2   8.999910E+1   -2.380000E+2   -2.380000E+2   -2.071049E-3   -1.432293E-5   -8.119080E-5   3.736901E-6   -3.738176E-6   -8.119074E-5   8.127675E-5   1.773648E+2   2.673639E+2   
2.924643E+3   2.039510E+1   2.039510E+1   -2.490000E+2   -2.490000E+2   8.999910E+1   -2.480000E+2   -2.480000E+2   -3.317276E-3   2.031441E-3   -8.389744E-5   3.114249E-6   -3.115567E-6   -8.389739E-5   8.395522E-5   1.778742E+2   2.678733E+2   
2.951501E+3   2.039410E+1   2.039410E+1   -2.590000E+2   -2.590000E+2   8.999910E+1   -2.580000E+2   -2.580000E+2   -4.415112E-3   3.319106E-3   -8.603658E-5   2.921673E-6   -2.923025E-6   -8.603654E-5   8.608617E-5   1.780551E+2   2.680542E+2   
2.978297E+3   2.041549E+1   2.041549E+1   -2.690000E+2   -2.690000E+2   8.999910E+1   -2.680000E+2   -2.680000E+2   -5.694244E-3   2.784050E-3   -8.717044E-5   4.136914E-6   -4.138283E-6   -8.717038E-5   8.726855E-5   1.772829E+2   2.672820E+2   
3.005097E+3   2.039999E+1   2.039999E+1   -2.790000E+2   -2.790000E+2   8.999910E+1   -2.780000E+2   -2.780000E+2   -7.040106E-3   4.821580E-3   -8.993849E-5   3.589265E-6   -3.590678E-6   -8.993843E-5   9.001008E-5   1.777147E+2   2.677138E+2   
3.031885E+3   2.040389E+1   2.040389E+1   -2.890000E+2   -2.890000E+2   8.999910E+1   -2.880000E+2   -2.880000E+2   -1.000911E-2   9.854927E-3   -9.564107E-5   2.062234E-6   -2.063736E-6   -9.564104E-5   9.566331E-5   1.787648E+2   2.687639E+2   
3.058697E+3   2.040121E+1   2.040121E+1   -2.990000E+2   -2.990000E+2   8.999910E+1   -2.980000E+2   -2.980000E+2   -9.776623E-3   7.149491E-3   -9.442488E-5   3.753814E-6   -3.755297E-6   -9.442482E-5   9.449947E-5   1.777234E+2   2.677225E+2   
3.085450E+3   2.039639E+1   2.039639E+1   -3.090000E+2   -3.090000E+2   8.999910E+1   -3.080000E+2   -3.080000E+2   -1.133456E-2   9.696790E-3   -9.764948E-5   2.994971E-6   -2.996505E-6   -9.764943E-5   9.769539E-5   1.782433E+2   2.682424E+2   
3.112296E+3   2.038369E+1   2.038369E+1   -3.190000E+2   -3.190000E+2   8.999910E+1   -3.180000E+2   -3.180000E+2   -1.316581E-2   1.031107E-2   -9.986205E-5   3.785436E-6   -3.787005E-6   -9.986199E-5   9.993377E-5   1.778291E+2   2.678282E+2   
3.139102E+3   2.038690E+1   2.038690E+1   -3.290000E+2   -3.290000E+2   8.999910E+1   -3.280000E+2   -3.280000E+2   -1.367223E-2   1.397723E-2   -1.030762E-4   1.509288E-6   -1.510907E-6   -1.030761E-4   1.030872E-4   1.791611E+2   2.691602E+2   
3.165907E+3   2.038180E+1   2.038180E+1   -3.390000E+2   -3.390000E+2   8.999910E+1   -3.380000E+2   -3.380000E+2   -1.488676E-2   1.312041E-2   -1.039681E-4   2.905947E-6   -2.907580E-6   -1.039680E-4   1.040087E-4   1.783990E+2   2.683981E+2   
3.192696E+3   2.038201E+1   2.038201E+1   -3.490000E+2   -3.490000E+2   8.999910E+1   -3.480000E+2   -3.480000E+2   -1.754466E-2   1.548977E-2   -1.078169E-4   3.036334E-6   -3.038027E-6   -1.078168E-4   1.078596E-4   1.783869E+2   2.683860E+2   
3.219501E+3   2.036541E+1   2.036541E+1   -3.590000E+2   -3.590000E+2   8.999910E+1   -3.580000E+2   -3.580000E+2   -1.863883E-2   1.694409E-2   -1.100566E-4   2.724005E-6   -2.725734E-6   -1.100565E-4   1.100903E-4   1.785822E+2   2.685813E+2   
3.246313E+3   2.036730E+1   2.036730E+1   -3.690000E+2   -3.690000E+2   8.999910E+1   -3.690000E+2   -3.690000E+2   -2.082811E-2   1.635817E-2   -1.118275E-4   4.602290E-6   -4.604047E-6   -1.118275E-4   1.119222E-4   1.776433E+2   2.676424E+2   
3.273107E+3   2.037179E+1   2.037179E+1   -3.790000E+2   -3.790000E+2   8.999910E+1   -3.780000E+2   -3.780000E+2   -2.072573E-2   1.735178E-2   -1.129228E-4   3.787748E-6   -3.789522E-6   -1.129228E-4   1.129863E-4   1.780789E+2   2.680780E+2   
3.299914E+3   2.035421E+1   2.035421E+1   -3.890000E+2   -3.890000E+2   8.999910E+1   -3.880000E+2   -3.880000E+2   -2.288302E-2   1.978543E-2   -1.164772E-4   3.525173E-6   -3.527003E-6   -1.164772E-4   1.165306E-4   1.782665E+2   2.682656E+2   
3.326708E+3   2.035931E+1   2.035931E+1   -3.990000E+2   -3.990000E+2   8.999910E+1   -3.980000E+2   -3.980000E+2   -2.256491E-2   2.008190E-2   -1.170588E-4   3.046095E-6   -3.047934E-6   -1.170588E-4   1.170985E-4   1.785094E+2   2.685085E+2   
3.353481E+3   2.035211E+1   2.035211E+1   -4.090000E+2   -4.090000E+2   8.999910E+1   -4.080000E+2   -4.080000E+2   -2.496688E-2   2.164653E-2   -1.202396E-4   3.564653E-6   -3.566542E-6   -1.202395E-4   1.202924E-4   1.783019E+2   2.683010E+2   
3.380289E+3   2.034649E+1   2.034649E+1   -4.190000E+2   -4.190000E+2   8.999910E+1   -4.180000E+2   -4.180000E+2   -2.644163E-2   2.350582E-2   -1.229835E-4   3.231887E-6   -3.233819E-6   -1.229835E-4   1.230260E-4   1.784947E+2   2.684938E+2   
3.407123E+3   2.036370E+1   2.036370E+1   -4.290000E+2   -4.290000E+2   8.999910E+1   -4.280000E+2   -4.280000E+2   -2.848282E-2   2.456313E-2   -1.256100E-4   3.856612E-6   -3.858585E-6   -1.256099E-4   1.256691E-4   1.782414E+2   2.682405E+2   
3.433904E+3   2.033999E+1   2.033999E+1   -4.390000E+2   -4.390000E+2   8.999910E+1   -4.380000E+2   -4.380000E+2   -2.972814E-2   2.589682E-2   -1.278760E-4   3.734120E-6   -3.736129E-6   -1.278759E-4   1.279305E-4   1.783274E+2   2.683265E+2   
3.460697E+3   2.034420E+1   2.034420E+1   -4.490000E+2   -4.490000E+2   8.999910E+1   -4.480000E+2   -4.480000E+2   -3.087380E-2   2.738435E-2   -1.301706E-4   3.434205E-6   -3.436250E-6   -1.301705E-4   1.302158E-4   1.784888E+2   2.684879E+2   
3.487509E+3   2.034219E+1   2.034219E+1   -4.590000E+2   -4.590000E+2   8.999910E+1   -4.580000E+2   -4.580000E+2   -3.261273E-2   2.887039E-2   -1.328602E-4   3.547451E-6   -3.549537E-6   -1.328601E-4   1.329075E-4   1.784705E+2   2.684696E+2   
3.514303E+3   2.034329E+1   2.034329E+1   -4.690000E+2   -4.690000E+2   8.999910E+1   -4.680000E+2   -4.680000E+2   -3.357283E-2   3.215200E-2   -1.361395E-4   1.856900E-6   -1.859039E-6   -1.361395E-4   1.361521E-4   1.792186E+2   2.692177E+2   
3.541102E+3   2.035269E+1   2.035269E+1   -4.790000E+2   -4.790000E+2   8.999910E+1   -4.780000E+2   -4.780000E+2   -3.526512E-2   2.451075E-2   -1.331581E-4   8.356775E-6   -8.358866E-6   -1.331579E-4   1.334200E-4   1.764089E+2   2.664080E+2   
3.567931E+3   2.035870E+1   2.035870E+1   -4.890000E+2   -4.890000E+2   8.999910E+1   -4.880000E+2   -4.880000E+2   -3.945961E-2   4.263976E-2   -1.477707E-4   -1.528870E-6   1.526549E-6   -1.477707E-4   1.477786E-4   -1.794072E+2   -8.940813E+1   
3.594704E+3   2.036450E+1   2.036450E+1   -4.990000E+2   -4.990000E+2   8.999910E+1   -4.980000E+2   -4.980000E+2   -3.818383E-2   2.456677E-2   -1.363622E-4   1.024565E-5   -1.024779E-5   -1.363621E-4   1.367466E-4   1.757031E+2   2.657022E+2   
3.621506E+3   2.036019E+1   2.036019E+1   -5.090000E+2   -5.090000E+2   8.999910E+1   -5.080000E+2   -5.080000E+2   -4.148282E-2   4.913487E-2   -1.543559E-4   -4.790521E-6   4.788096E-6   -1.543560E-4   1.544303E-4   -1.782224E+2   -8.822326E+1   
3.648301E+3   2.037249E+1   2.037249E+1   -5.190000E+2   -5.190000E+2   8.999910E+1   -5.180000E+2   -5.180000E+2   -3.771643E-2   3.434097E-2   -1.433114E-4   2.947795E-6   -2.950046E-6   -1.433113E-4   1.433417E-4   1.788216E+2   2.688207E+2   
3.675128E+3   2.036721E+1   2.036721E+1   -5.290000E+2   -5.290000E+2   8.999910E+1   -5.280000E+2   -5.280000E+2   -4.274764E-2   3.708209E-2   -1.489739E-4   4.465340E-6   -4.467680E-6   -1.489739E-4   1.490409E-4   1.782831E+2   2.682822E+2   
3.701907E+3   2.038641E+1   2.038641E+1   -5.390000E+2   -5.390000E+2   8.999910E+1   -5.380000E+2   -5.380000E+2   -4.477908E-2   3.377788E-2   -1.488988E-4   8.150659E-6   -8.152998E-6   -1.488987E-4   1.491217E-4   1.768668E+2   2.668659E+2   
3.728693E+3   2.038171E+1   2.038171E+1   -5.490000E+2   -5.490000E+2   8.999910E+1   -5.490000E+2   -5.490000E+2   -4.642389E-2   4.161239E-2   -1.555095E-4   3.728824E-6   -3.731267E-6   -1.555095E-4   1.555542E-4   1.786264E+2   2.686255E+2   
3.755542E+3   2.038070E+1   2.038070E+1   -5.590000E+2   -5.590000E+2   8.999910E+1   -5.580000E+2   -5.580000E+2   -4.935087E-2   4.608173E-2   -1.607745E-4   2.574209E-6   -2.576734E-6   -1.607745E-4   1.607951E-4   1.790827E+2   2.690818E+2   
3.782456E+3   2.036111E+1   2.036111E+1   -5.690000E+2   -5.690000E+2   8.999910E+1   -5.690000E+2   -5.690000E+2   -4.844194E-2   4.478400E-2   -1.600377E-4   2.800938E-6   -2.803452E-6   -1.600377E-4   1.600622E-4   1.789973E+2   2.689964E+2   
3.809259E+3   2.035751E+1   2.035751E+1   -5.790000E+2   -5.790000E+2   8.999910E+1   -5.780000E+2   -5.780000E+2   -5.092680E-2   4.514537E-2   -1.624692E-4   4.228259E-6   -4.230811E-6   -1.624691E-4   1.625242E-4   1.785092E+2   2.685083E+2   
3.836033E+3   2.035839E+1   2.035839E+1   -5.890000E+2   -5.890000E+2   8.999910E+1   -5.890000E+2   -5.890000E+2   -5.191311E-2   4.488057E-2   -1.636357E-4   5.045066E-6   -5.047637E-6   -1.636356E-4   1.637134E-4   1.782341E+2   2.682332E+2   
3.862846E+3   2.037219E+1   2.037219E+1   -5.990000E+2   -5.990000E+2   8.999910E+1   -5.980000E+2   -5.980000E+2   -5.316911E-2   4.671032E-2   -1.661543E-4   4.586079E-6   -4.588689E-6   -1.661542E-4   1.662176E-4   1.784190E+2   2.684181E+2   
3.889649E+3   2.036419E+1   2.036419E+1   -6.090000E+2   -6.090000E+2   8.999910E+1   -6.080000E+2   -6.080000E+2   -5.596167E-2   4.842484E-2   -1.696883E-4   5.270538E-6   -5.273203E-6   -1.696883E-4   1.697702E-4   1.782210E+2   2.682201E+2   
3.916451E+3   2.036309E+1   2.036309E+1   -6.190000E+2   -6.190000E+2   8.999910E+1   -6.190000E+2   -6.190000E+2   -5.732733E-2   5.160563E-2   -1.732371E-4   3.927655E-6   -3.930376E-6   -1.732371E-4   1.732816E-4   1.787012E+2   2.687003E+2   
3.943254E+3   2.037011E+1   2.037011E+1   -6.290000E+2   -6.290000E+2   8.999910E+1   -6.290000E+2   -6.290000E+2   -5.835509E-2   5.403713E-2   -1.760363E-4   2.881968E-6   -2.884733E-6   -1.760363E-4   1.760599E-4   1.790621E+2   2.690612E+2   
3.970049E+3   2.036001E+1   2.036001E+1   -6.390000E+2   -6.390000E+2   8.999910E+1   -6.380000E+2   -6.380000E+2   -6.015098E-2   5.416328E-2   -1.778626E-4   3.996118E-6   -3.998912E-6   -1.778625E-4   1.779074E-4   1.787129E+2   2.687120E+2   
3.996851E+3   2.034130E+1   2.034130E+1   -6.490000E+2   -6.490000E+2   8.999910E+1   -6.490000E+2   -6.490000E+2   -6.315472E-2   5.489304E-2   -1.809901E-4   5.514885E-6   -5.517727E-6   -1.809901E-4   1.810741E-4   1.782547E+2   2.682538E+2   
4.023653E+3   2.033120E+1   2.033120E+1   -6.600000E+2   -6.600000E+2   8.999910E+1   -6.590000E+2   -6.590000E+2   -6.438782E-2   5.729712E-2   -1.839094E-4   4.631114E-6   -4.634003E-6   -1.839094E-4   1.839677E-4   1.785575E+2   2.685566E+2   
4.050455E+3   2.032769E+1   2.032769E+1   -6.690000E+2   -6.690000E+2   8.999910E+1   -6.690000E+2   -6.690000E+2   -6.552861E-2   5.701497E-2   -1.851072E-4   5.572392E-6   -5.575299E-6   -1.851071E-4   1.851911E-4   1.782757E+2   2.682748E+2   
4.077245E+3   2.034011E+1   2.034011E+1   -6.790000E+2   -6.790000E+2   8.999910E+1   -6.790000E+2   -6.790000E+2   -6.663437E-2   5.937034E-2   -1.879114E-4   4.634430E-6   -4.637381E-6   -1.879113E-4   1.879685E-4   1.785872E+2   2.685863E+2   
4.104053E+3   2.033129E+1   2.033129E+1   -6.890000E+2   -6.890000E+2   8.999910E+1   -6.890000E+2   -6.890000E+2   -6.726813E-2   6.237192E-2   -1.907999E-4   2.914123E-6   -2.917120E-6   -1.907998E-4   1.908221E-4   1.791250E+2   2.691241E+2   
4.130847E+3   2.033590E+1   2.033590E+1   -6.990000E+2   -6.990000E+2   8.999910E+1   -6.990000E+2   -6.990000E+2   -7.103819E-2   6.318120E-2   -1.944270E-4   4.914236E-6   -4.917290E-6   -1.944269E-4   1.944891E-4   1.785521E+2   2.685512E+2   
4.157640E+3   2.033480E+1   2.033480E+1   -7.100000E+2   -7.100000E+2   8.999910E+1   -7.090000E+2   -7.090000E+2   -7.323567E-2   6.488873E-2   -1.975595E-4   5.190244E-6   -5.193347E-6   -1.975595E-4   1.976277E-4   1.784951E+2   2.684942E+2   
4.184416E+3   2.034481E+1   2.034481E+1   -7.190000E+2   -7.190000E+2   8.999910E+1   -7.190000E+2   -7.190000E+2   -7.318692E-2   6.592228E-2   -1.987764E-4   4.379907E-6   -4.383029E-6   -1.987763E-4   1.988246E-4   1.787377E+2   2.687368E+2   
4.211257E+3   2.035510E+1   2.035510E+1   -7.290000E+2   -7.290000E+2   8.999910E+1   -7.290000E+2   -7.290000E+2   -7.591487E-2   6.884556E-2   -2.030142E-4   4.169392E-6   -4.172581E-6   -2.030142E-4   2.030570E-4   1.788235E+2   2.688226E+2   
4.238056E+3   2.034741E+1   2.034741E+1   -7.400000E+2   -7.400000E+2   8.999910E+1   -7.390000E+2   -7.390000E+2   -7.668913E-2   7.128102E-2   -2.056466E-4   2.944828E-6   -2.948059E-6   -2.056466E-4   2.056677E-4   1.791796E+2   2.691787E+2   
4.264860E+3   2.034420E+1   2.034420E+1   -7.500000E+2   -7.500000E+2   8.999910E+1   -7.490000E+2   -7.490000E+2   -7.984520E-2   7.258179E-2   -2.091677E-4   4.172784E-6   -4.176070E-6   -2.091676E-4   2.092093E-4   1.788571E+2   2.688562E+2   
4.291645E+3   2.035510E+1   2.035510E+1   -7.600000E+2   -7.600000E+2   8.999910E+1   -7.590000E+2   -7.590000E+2   -8.255062E-2   7.435788E-2   -2.126816E-4   4.753415E-6   -4.756755E-6   -2.126815E-4   2.127347E-4   1.787197E+2   2.687188E+2   
4.318450E+3   2.035659E+1   2.035659E+1   -7.690000E+2   -7.690000E+2   8.999910E+1   -7.690000E+2   -7.690000E+2   -8.457660E-2   7.643045E-2   -2.159252E-4   4.653559E-6   -4.656951E-6   -2.159252E-4   2.159754E-4   1.787654E+2   2.687645E+2   
4.345254E+3   2.034789E+1   2.034789E+1   -7.800000E+2   -7.800000E+2   8.999910E+1   -7.790000E+2   -7.790000E+2   -8.551474E-2   8.039979E-2   -2.196149E-4   2.464095E-6   -2.467544E-6   -2.196148E-4   2.196287E-4   1.793572E+2   2.693563E+2   
4.372055E+3   2.037341E+1   2.037341E+1   -7.900000E+2   -7.900000E+2   8.999910E+1   -7.890000E+2   -7.890000E+2   -8.916237E-2   8.043730E-2   -2.226834E-4   4.921929E-6   -4.925427E-6   -2.226833E-4   2.227378E-4   1.787338E+2   2.687329E+2   
4.398880E+3   2.039791E+1   2.039791E+1   -7.990000E+2   -7.990000E+2   8.999910E+1   -7.990000E+2   -7.990000E+2   -8.905024E-2   8.230965E-2   -2.243762E-4   3.477656E-6   -3.481181E-6   -2.243762E-4   2.244032E-4   1.791120E+2   2.691111E+2   
4.425648E+3   2.037731E+1   2.037731E+1   -8.090000E+2   -8.090000E+2   8.999910E+1   -8.090000E+2   -8.090000E+2   -8.947740E-2   8.166034E-2   -2.248708E-4   4.181432E-6   -4.184964E-6   -2.248708E-4   2.249097E-4   1.789347E+2   2.689338E+2   
4.452457E+3   2.036831E+1   2.036831E+1   -8.190000E+2   -8.190000E+2   8.999910E+1   -8.190000E+2   -8.190000E+2   -9.206709E-2   8.460073E-2   -2.290270E-4   3.862840E-6   -3.866438E-6   -2.290269E-4   2.290595E-4   1.790337E+2   2.690328E+2   
4.479259E+3   2.036279E+1   2.036279E+1   -8.290000E+2   -8.290000E+2   8.999910E+1   -8.290000E+2   -8.290000E+2   -9.415436E-2   8.528386E-2   -2.314529E-4   4.782726E-6   -4.786362E-6   -2.314529E-4   2.315024E-4   1.788162E+2   2.688153E+2   
4.506069E+3   2.034210E+1   2.034210E+1   -8.390000E+2   -8.390000E+2   8.999910E+1   -8.390000E+2   -8.390000E+2   -9.501425E-2   8.749840E-2   -2.340060E-4   3.773013E-6   -3.776689E-6   -2.340059E-4   2.340364E-4   1.790763E+2   2.690754E+2   
4.532811E+3   2.037130E+1   2.037130E+1   -8.500000E+2   -8.500000E+2   8.999910E+1   -8.490000E+2   -8.490000E+2   -9.802168E-2   8.949085E-2   -2.378552E-4   4.411277E-6   -4.415013E-6   -2.378551E-4   2.378961E-4   1.789375E+2   2.689366E+2   
4.559661E+3   2.035021E+1   2.035021E+1   -8.590000E+2   -8.590000E+2   8.999910E+1   -8.580000E+2   -8.580000E+2   -1.003761E-1   9.539326E-2   -2.436236E-4   1.851124E-6   -1.854951E-6   -2.436235E-4   2.436306E-4   1.795647E+2   2.695638E+2   
4.586476E+3   2.035909E+1   2.035909E+1   -8.690000E+2   -8.690000E+2   8.999910E+1   -8.690000E+2   -8.690000E+2   -1.017421E-1   8.891585E-2   -2.412046E-4   7.300875E-6   -7.304664E-6   -2.412045E-4   2.413151E-4   1.782663E+2   2.682654E+2   
4.613225E+3   2.035589E+1   2.035589E+1   -8.790000E+2   -8.790000E+2   8.999910E+1   -8.790000E+2   -8.790000E+2   -1.057925E-1   9.621348E-2   -2.490281E-4   4.932594E-6   -4.936506E-6   -2.490280E-4   2.490769E-4   1.788653E+2   2.688644E+2   
4.640072E+3   2.035360E+1   2.035360E+1   -8.890000E+2   -8.890000E+2   8.999910E+1   -8.880000E+2   -8.880000E+2   -1.068824E-1   1.024480E-1   -2.541576E-4   1.260423E-6   -1.264416E-6   -2.541576E-4   2.541607E-4   1.797159E+2   2.697150E+2   
4.666887E+3   2.034179E+1   2.034179E+1   -8.990000E+2   -8.990000E+2   8.999910E+1   -8.990000E+2   -8.990000E+2   -1.106866E-1   1.064619E-1   -2.598487E-4   1.025575E-6   -1.029657E-6   -2.598487E-4   2.598507E-4   1.797739E+2   2.697730E+2   
4.693641E+3   2.034979E+1   2.034979E+1   -9.090000E+2   -9.090000E+2   8.999910E+1   -9.090000E+2   -9.090000E+2   -1.135373E-1   1.073233E-1   -2.628945E-4   2.350453E-6   -2.354582E-6   -2.628944E-4   2.629050E-4   1.794878E+2   2.694869E+2   
4.720455E+3   2.036361E+1   2.036361E+1   -9.190000E+2   -9.190000E+2   8.999910E+1   -9.190000E+2   -9.190000E+2   -1.169557E-1   1.068903E-1   -2.655193E-4   4.979934E-6   -4.984105E-6   -2.655192E-4   2.655660E-4   1.789255E+2   2.689246E+2   
4.747282E+3   2.035739E+1   2.035739E+1   -9.290000E+2   -9.290000E+2   8.999910E+1   -9.290000E+2   -9.290000E+2   -1.188159E-1   1.106390E-1   -2.696880E-4   3.586118E-6   -3.590354E-6   -2.696879E-4   2.697118E-4   1.792382E+2   2.692373E+2   
4.774070E+3   2.034771E+1   2.034771E+1   -9.390000E+2   -9.390000E+2   8.999910E+1   -9.390000E+2   -9.390000E+2   -1.213145E-1   1.133426E-1   -2.736370E-4   3.370719E-6   -3.375017E-6   -2.736369E-4   2.736577E-4   1.792943E+2   2.692934E+2   
4.800873E+3   2.035201E+1   2.035201E+1   -9.490000E+2   -9.490000E+2   8.999910E+1   -9.490000E+2   -9.490000E+2   -1.252539E-1   1.178845E-1   -2.796836E-4   2.863486E-6   -2.867879E-6   -2.796835E-4   2.796982E-4   1.794134E+2   2.694125E+2   
4.827662E+3   2.036569E+1   2.036569E+1   -9.590000E+2   -9.590000E+2   8.999910E+1   -9.590000E+2   -9.590000E+2   -1.269685E-1   1.230534E-1   -2.846326E-4   3.697086E-7   -3.741796E-7   -2.846326E-4   2.846329E-4   1.799256E+2   2.699247E+2   
4.854484E+3   2.035781E+1   2.035781E+1   -9.690000E+2   -9.690000E+2   8.999910E+1   -9.690000E+2   -9.690000E+2   -1.293896E-1   1.257747E-1   -2.885409E-4   8.812067E-8   -9.265306E-8   -2.885409E-4   2.885409E-4   1.799825E+2   2.699816E+2   
4.881262E+3   2.037750E+1   2.037750E+1   -9.800000E+2   -9.800000E+2   8.999910E+1   -9.790000E+2   -9.790000E+2   -1.339549E-1   1.302775E-1   -2.949811E-4   4.306175E-8   -4.769530E-8   -2.949811E-4   2.949811E-4   1.799916E+2   2.699907E+2   
4.908085E+3   2.037231E+1   2.037231E+1   -9.890000E+2   -9.890000E+2   8.999910E+1   -9.880000E+2   -9.880000E+2   -1.379047E-1   1.314487E-1   -2.988908E-4   1.918430E-6   -1.923125E-6   -2.988908E-4   2.988970E-4   1.796323E+2   2.696314E+2   
4.934890E+3   2.037670E+1   2.037670E+1   -9.990000E+2   -9.990000E+2   8.999910E+1   -9.980000E+2   -9.980000E+2   -1.414011E-1   1.385025E-1   -3.061939E-4   -6.631625E-7   6.583528E-7   -3.061939E-4   3.061946E-4   -1.798759E+2   -8.987681E+1   
4.961794E+3   2.036709E+1   2.036709E+1   -1.009000E+3   -1.009000E+3   8.999910E+1   -1.009000E+3   -1.009000E+3   -1.463266E-1   1.419847E-1   -3.123049E-4   2.548474E-7   -2.597530E-7   -3.123048E-4   3.123050E-4   1.799532E+2   2.699523E+2   
4.988752E+3   2.036221E+1   2.036221E+1   -1.019000E+3   -1.019000E+3   8.999910E+1   -1.018000E+3   -1.018000E+3   -1.499208E-1   1.461526E-1   -3.178290E-4   -2.243043E-7   2.193118E-7   -3.178290E-4   3.178290E-4   -1.799596E+2   -8.996046E+1   
5.015695E+3   2.035009E+1   2.035009E+1   -1.029000E+3   -1.029000E+3   8.999910E+1   -1.028000E+3   -1.028000E+3   -1.537649E-1   1.520811E-1   -3.246688E-4   -1.773004E-6   1.767904E-6   -3.246688E-4   3.246736E-4   -1.796871E+2   -8.968801E+1   
5.042640E+3   2.034081E+1   2.034081E+1   -1.039000E+3   -1.039000E+3   8.999910E+1   -1.038000E+3   -1.038000E+3   -1.587586E-1   1.568878E-1   -3.315826E-4   -1.734144E-6   1.728936E-6   -3.315827E-4   3.315872E-4   -1.797004E+2   -8.970125E+1   
5.069555E+3   2.034799E+1   2.034799E+1   -1.049000E+3   -1.049000E+3   8.999910E+1   -1.048000E+3   -1.048000E+3   -1.642313E-1   1.637450E-1   -3.400834E-4   -2.804707E-6   2.799365E-6   -3.400834E-4   3.400949E-4   -1.795275E+2   -8.952839E+1   
5.096474E+3   2.035180E+1   2.035180E+1   -1.059000E+3   -1.059000E+3   8.999910E+1   -1.059000E+3   -1.059000E+3   -1.698463E-1   1.677927E-1   -3.470040E-4   -1.805476E-6   1.800025E-6   -3.470041E-4   3.470087E-4   -1.797019E+2   -8.970279E+1   
5.123415E+3   2.034881E+1   2.034881E+1   -1.069000E+3   -1.069000E+3   8.999910E+1   -1.068000E+3   -1.068000E+3   -1.730832E-1   1.775176E-1   -3.557233E-4   -6.440911E-6   6.435323E-6   -3.557234E-4   3.557816E-4   -1.789627E+2   -8.896359E+1   
5.150348E+3   2.033779E+1   2.033779E+1   -1.079000E+3   -1.079000E+3   8.999910E+1   -1.078000E+3   -1.078000E+3   -1.778911E-1   1.807599E-1   -3.615466E-4   -5.430958E-6   5.425279E-6   -3.615467E-4   3.615874E-4   -1.791394E+2   -8.914030E+1   
5.177305E+3   2.031970E+1   2.031970E+1   -1.089000E+3   -1.089000E+3   8.999910E+1   -1.088000E+3   -1.088000E+3   -1.836257E-1   1.855955E-1   -3.689729E-4   -4.897847E-6   4.892052E-6   -3.689729E-4   3.690054E-4   -1.792395E+2   -8.924038E+1   
5.204242E+3   2.033419E+1   2.033419E+1   -1.099000E+3   -1.099000E+3   8.999910E+1   -1.099000E+3   -1.099000E+3   -1.880646E-1   1.933348E-1   -3.773897E-4   -7.311728E-6   7.305799E-6   -3.773898E-4   3.774605E-4   -1.788901E+2   -8.889096E+1   
5.231181E+3   2.032931E+1   2.032931E+1   -1.109000E+3   -1.109000E+3   8.999910E+1   -1.108000E+3   -1.108000E+3   -1.926831E-1   1.995060E-1   -3.848353E-4   -8.488291E-6   8.482246E-6   -3.848354E-4   3.849289E-4   -1.787364E+2   -8.873733E+1   
5.258220E+3   2.032501E+1   2.032501E+1   -1.119000E+3   -1.119000E+3   8.999910E+1   -1.118000E+3   -1.118000E+3   -1.980603E-1   2.036229E-1   -3.915789E-4   -7.697905E-6   7.691754E-6   -3.915790E-4   3.916545E-4   -1.788738E+2   -8.887469E+1   
5.285207E+3   2.031429E+1   2.031429E+1   -1.129000E+3   -1.129000E+3   8.999910E+1   -1.128000E+3   -1.128000E+3   -2.020967E-1   2.091096E-1   -3.982740E-4   -8.802340E-6   8.796084E-6   -3.982742E-4   3.983713E-4   -1.787339E+2   -8.873480E+1   
5.312225E+3   2.032260E+1   2.032260E+1   -1.139000E+3   -1.139000E+3   8.999910E+1   -1.138000E+3   -1.138000E+3   -2.039410E-1   2.144549E-1   -4.034187E-4   -1.133002E-5   1.132368E-5   -4.034189E-4   4.035778E-4   -1.783913E+2   -8.839217E+1   
5.339175E+3   2.032629E+1   2.032629E+1   -1.149000E+3   -1.149000E+3   8.999910E+1   -1.148000E+3   -1.148000E+3   -2.069109E-1   2.146274E-1   -4.061183E-4   -9.437895E-6   9.431516E-6   -4.061184E-4   4.062279E-4   -1.786687E+2   -8.866963E+1   
5.366132E+3   2.032061E+1   2.032061E+1   -1.159000E+3   -1.159000E+3   8.999910E+1   -1.158000E+3   -1.158000E+3   -2.076775E-1   2.164163E-1   -4.083461E-4   -1.021305E-5   1.020663E-5   -4.083463E-4   4.084738E-4   -1.785673E+2   -8.856819E+1   
5.393171E+3   2.029781E+1   2.029781E+1   -1.169000E+3   -1.169000E+3   8.999910E+1   -1.169000E+3   -1.169000E+3   -2.078786E-1   2.165400E-1   -4.092286E-4   -1.021489E-5   1.020846E-5   -4.092287E-4   4.093560E-4   -1.785701E+2   -8.857102E+1   
5.420137E+3   2.031851E+1   2.031851E+1   -1.179000E+3   -1.179000E+3   8.999910E+1   -1.179000E+3   -1.179000E+3   -2.085800E-1   2.156640E-1   -4.097661E-4   -9.161175E-6   9.154739E-6   -4.097663E-4   4.098685E-4   -1.787192E+2   -8.872015E+1   
5.447151E+3   2.031429E+1   2.031429E+1   -1.189000E+3   -1.189000E+3   8.999910E+1   -1.189000E+3   -1.189000E+3   -2.083561E-1   2.165638E-1   -4.107834E-4   -9.999143E-6   9.992691E-6   -4.107835E-4   4.109050E-4   -1.786056E+2   -8.860650E+1   
5.474131E+3   2.032351E+1   2.032351E+1   -1.199000E+3   -1.199000E+3   8.999910E+1   -1.198000E+3   -1.198000E+3   -2.067058E-1   2.150165E-1   -4.092755E-4   -1.010196E-5   1.009553E-5   -4.092756E-4   4.094001E-4   -1.785861E+2   -8.858698E+1   
5.501154E+3   2.031909E+1   2.031909E+1   -1.209000E+3   -1.209000E+3   8.999910E+1   -1.208000E+3   -1.208000E+3   -2.057710E-1   2.134162E-1   -4.082734E-4   -9.675493E-6   9.669080E-6   -4.082735E-4   4.083880E-4   -1.786424E+2   -8.864333E+1   
5.528106E+3   2.033569E+1   2.033569E+1   -1.219000E+3   -1.219000E+3   8.999910E+1   -1.218000E+3   -1.218000E+3   -2.064304E-1   2.147343E-1   -4.101387E-4   -1.019407E-5   1.018763E-5   -4.101389E-4   4.102654E-4   -1.785762E+2   -8.857710E+1   
5.555059E+3   2.032211E+1   2.032211E+1   -1.229000E+3   -1.229000E+3   8.999910E+1   -1.228000E+3   -1.228000E+3   -2.062497E-1   2.148925E-1   -4.107266E-4   -1.048040E-5   1.047395E-5   -4.107267E-4   4.108603E-4   -1.785383E+2   -8.853922E+1   
5.582002E+3   2.032891E+1   2.032891E+1   -1.239000E+3   -1.239000E+3   8.999910E+1   -1.238000E+3   -1.238000E+3   -2.076282E-1   2.142950E-1   -4.118881E-4   -9.152242E-6   9.145772E-6   -4.118883E-4   4.119898E-4   -1.787271E+2   -8.872799E+1   
5.609022E+3   2.032430E+1   2.032430E+1   -1.249000E+3   -1.249000E+3   8.999910E+1   -1.248000E+3   -1.248000E+3   -2.062528E-1   2.131786E-1   -4.108910E-4   -9.372105E-6   9.365651E-6   -4.108911E-4   4.109978E-4   -1.786934E+2   -8.869425E+1   
5.636005E+3   2.033749E+1   2.033749E+1   -1.259000E+3   -1.259000E+3   8.999910E+1   -1.258000E+3   -1.258000E+3   -2.058186E-1   2.127078E-1   -4.109210E-4   -9.392255E-6   9.385801E-6   -4.109211E-4   4.110283E-4   -1.786906E+2   -8.869154E+1   
5.663028E+3   2.032281E+1   2.032281E+1   -1.269000E+3   -1.269000E+3   8.999910E+1   -1.268000E+3   -1.268000E+3   -2.052588E-1   2.142331E-1   -4.121006E-4   -1.090338E-5   1.089691E-5   -4.121008E-4   4.122449E-4   -1.784844E+2   -8.848532E+1   
5.690004E+3   2.032101E+1   2.032101E+1   -1.279000E+3   -1.279000E+3   8.999910E+1   -1.278000E+3   -1.278000E+3   -2.049959E-1   2.136624E-1   -4.121832E-4   -1.073429E-5   1.072781E-5   -4.121834E-4   4.123230E-4   -1.785082E+2   -8.850911E+1   
5.717015E+3   2.032198E+1   2.032198E+1   -1.289000E+3   -1.289000E+3   8.999910E+1   -1.289000E+3   -1.289000E+3   -2.041845E-1   2.127563E-1   -4.117535E-4   -1.071520E-5   1.070873E-5   -4.117537E-4   4.118929E-4   -1.785093E+2   -8.851021E+1   
5.744011E+3   2.033361E+1   2.033361E+1   -1.299000E+3   -1.299000E+3   8.999910E+1   -1.298000E+3   -1.298000E+3   -2.042259E-1   2.118708E-1   -4.117836E-4   -1.010835E-5   1.010189E-5   -4.117838E-4   4.119077E-4   -1.785938E+2   -8.859470E+1   
5.771017E+3   2.033318E+1   2.033318E+1   -1.309000E+3   -1.309000E+3   8.999910E+1   -1.308000E+3   -1.308000E+3   -2.040224E-1   2.119939E-1   -4.123346E-4   -1.038589E-5   1.037942E-5   -4.123347E-4   4.124654E-4   -1.785571E+2   -8.855804E+1   
5.797986E+3   2.033801E+1   2.033801E+1   -1.319000E+3   -1.319000E+3   8.999910E+1   -1.318000E+3   -1.318000E+3   -2.036122E-1   2.114582E-1   -4.123406E-4   -1.034366E-5   1.033719E-5   -4.123407E-4   4.124703E-4   -1.785630E+2   -8.856392E+1   
5.824925E+3   2.031310E+1   2.031310E+1   -1.329000E+3   -1.329000E+3   8.999910E+1   -1.329000E+3   -1.329000E+3   -2.039401E-1   2.107233E-1   -4.127771E-4   -9.653632E-6   9.647148E-6   -4.127772E-4   4.128899E-4   -1.786603E+2   -8.866117E+1   
5.851877E+3   2.032031E+1   2.032031E+1   -1.339000E+3   -1.339000E+3   8.999910E+1   -1.338000E+3   -1.338000E+3   -2.038435E-1   2.118784E-1   -4.139760E-4   -1.057771E-5   1.057121E-5   -4.139762E-4   4.141111E-4   -1.785363E+2   -8.853722E+1   
5.878917E+3   2.033581E+1   2.033581E+1   -1.349000E+3   -1.349000E+3   8.999910E+1   -1.349000E+3   -1.349000E+3   -2.020872E-1   2.116718E-1   -4.133479E-4   -1.170699E-5   1.170049E-5   -4.133481E-4   4.135137E-4   -1.783777E+2   -8.837858E+1   
5.905864E+3   2.032620E+1   2.032620E+1   -1.359000E+3   -1.359000E+3   8.999910E+1   -1.358000E+3   -1.358000E+3   -2.028285E-1   2.103043E-1   -4.135474E-4   -1.027493E-5   1.026844E-5   -4.135475E-4   4.136750E-4   -1.785767E+2   -8.857763E+1   
5.932765E+3   2.033129E+1   2.033129E+1   -1.369000E+3   -1.369000E+3   8.999910E+1   -1.368000E+3   -1.368000E+3   -2.029757E-1   2.117383E-1   -4.151424E-4   -1.123075E-5   1.122423E-5   -4.151425E-4   4.152942E-4   -1.784504E+2   -8.845127E+1   
5.959712E+3   2.032491E+1   2.032491E+1   -1.379000E+3   -1.379000E+3   8.999910E+1   -1.378000E+3   -1.378000E+3   -2.028578E-1   2.109055E-1   -4.151598E-4   -1.077659E-5   1.077007E-5   -4.151600E-4   4.152996E-4   -1.785131E+2   -8.851397E+1   
5.986662E+3   2.033059E+1   2.033059E+1   -1.389000E+3   -1.389000E+3   8.999910E+1   -1.388000E+3   -1.388000E+3   -2.012084E-1   2.092315E-1   -4.136352E-4   -1.079464E-5   1.078814E-5   -4.136354E-4   4.137761E-4   -1.785051E+2   -8.850599E+1   
6.013598E+3   2.034039E+1   2.034039E+1   -1.399000E+3   -1.399000E+3   8.999910E+1   -1.398000E+3   -1.398000E+3   -2.033334E-1   2.105597E-1   -4.164850E-4   -1.030218E-5   1.029564E-5   -4.164852E-4   4.166124E-4   -1.785830E+2   -8.858392E+1   
6.040541E+3   2.034631E+1   2.034631E+1   -1.409000E+3   -1.409000E+3   8.999910E+1   -1.408000E+3   -1.408000E+3   -2.011052E-1   2.110237E-1   -4.158952E-4   -1.222600E-5   1.221947E-5   -4.158954E-4   4.160749E-4   -1.783162E+2   -8.831707E+1   
6.067486E+3   2.034438E+1   2.034438E+1   -1.419000E+3   -1.419000E+3   8.999910E+1   -1.418000E+3   -1.418000E+3   -2.025178E-1   2.090127E-1   -4.162061E-4   -9.880044E-6   9.873506E-6   -4.162063E-4   4.163234E-4   -1.786401E+2   -8.864105E+1   
6.094423E+3   2.034219E+1   2.034219E+1   -1.429000E+3   -1.429000E+3   8.999910E+1   -1.428000E+3   -1.428000E+3   -2.009929E-1   2.109463E-1   -4.169940E-4   -1.234873E-5   1.234218E-5   -4.169941E-4   4.171768E-4   -1.783038E+2   -8.830466E+1   
6.121427E+3   2.034579E+1   2.034579E+1   -1.439000E+3   -1.439000E+3   8.999910E+1   -1.438000E+3   -1.438000E+3   -2.014631E-1   2.072927E-1   -4.156608E-4   -9.502166E-6   9.495637E-6   -4.156610E-4   4.157694E-4   -1.786904E+2   -8.869132E+1   
6.148403E+3   2.035061E+1   2.035061E+1   -1.449000E+3   -1.449000E+3   8.999910E+1   -1.448000E+3   -1.448000E+3   -2.009833E-1   2.096075E-1   -4.173816E-4   -1.151307E-5   1.150651E-5   -4.173818E-4   4.175404E-4   -1.784200E+2   -8.842085E+1   
6.175360E+3   2.035781E+1   2.035781E+1   -1.459000E+3   -1.459000E+3   8.999910E+1   -1.458000E+3   -1.458000E+3   -2.004079E-1   2.091925E-1   -4.173519E-4   -1.167043E-5   1.166388E-5   -4.173521E-4   4.175150E-4   -1.783983E+2   -8.839915E+1   
6.202387E+3   2.036410E+1   2.036410E+1   -1.469000E+3   -1.469000E+3   8.999910E+1   -1.468000E+3   -1.468000E+3   -2.027295E-1   2.078530E-1   -4.186845E-4   -9.165357E-6   9.158780E-6   -4.186846E-4   4.187848E-4   -1.787459E+2   -8.874685E+1   
6.230046E+3   2.035281E+1   2.035281E+1   -1.479000E+3   -1.479000E+3   8.999910E+1   -1.478000E+3   -1.478000E+3   -1.994652E-1   2.068219E-1   -4.164793E-4   -1.075735E-5   1.075080E-5   -4.164795E-4   4.166182E-4   -1.785204E+2   -8.852132E+1   
6.257088E+3   2.034420E+1   2.034420E+1   -1.489000E+3   -1.489000E+3   8.999910E+1   -1.488000E+3   -1.488000E+3   -2.002269E-1   2.093671E-1   -4.191711E-4   -1.206777E-5   1.206119E-5   -4.191713E-4   4.193448E-4   -1.783509E+2   -8.835183E+1   
6.284096E+3   2.033160E+1   2.033160E+1   -1.499000E+3   -1.499000E+3   8.999910E+1   -1.498000E+3   -1.498000E+3   -1.999128E-1   2.083521E-1   -4.189451E-4   -1.162177E-5   1.161519E-5   -4.189452E-4   4.191062E-4   -1.784110E+2   -8.841189E+1   
6.311042E+3   2.033071E+1   2.033071E+1   -1.509000E+3   -1.509000E+3   8.999910E+1   -1.508000E+3   -1.508000E+3   -2.006109E-1   2.107029E-1   -4.214743E-4   -1.283971E-5   1.283309E-5   -4.214745E-4   4.216698E-4   -1.782551E+2   -8.825599E+1   
6.338482E+3   2.034899E+1   2.034899E+1   -1.518000E+3   -1.518000E+3   8.999910E+1   -1.518000E+3   -1.518000E+3   -1.964254E-1   2.065346E-1   -4.167157E-4   -1.286528E-5   1.285873E-5   -4.167159E-4   4.169142E-4   -1.782317E+2   -8.823257E+1   
6.365473E+3   2.034600E+1   2.034600E+1   -1.529000E+3   -1.529000E+3   8.999910E+1   -1.528000E+3   -1.528000E+3   -1.954515E-1   1.941377E-1   -4.090162E-4   -4.872921E-6   4.866496E-6   -4.090163E-4   4.090452E-4   -1.793174E+2   -8.931832E+1   
6.393213E+3   2.033859E+1   2.033859E+1   -1.538000E+3   -1.538000E+3   8.999910E+1   -1.537000E+3   -1.537000E+3   -1.963943E-1   2.038349E-1   -4.161871E-4   -1.108246E-5   1.107593E-5   -4.161873E-4   4.163347E-4   -1.784747E+2   -8.847556E+1   
6.420147E+3   2.034051E+1   2.034051E+1   -1.549000E+3   -1.549000E+3   8.999910E+1   -1.548000E+3   -1.548000E+3   -1.962231E-1   2.022871E-1   -4.157882E-4   -1.016739E-5   1.016086E-5   -4.157884E-4   4.159125E-4   -1.785992E+2   -8.860011E+1   
6.447685E+3   2.032211E+1   2.032211E+1   -1.558000E+3   -1.558000E+3   8.999910E+1   -1.558000E+3   -1.558000E+3   -1.967222E-1   2.059712E-1   -4.190086E-4   -1.246127E-5   1.245468E-5   -4.190088E-4   4.191938E-4   -1.782965E+2   -8.829743E+1   
6.474688E+3   2.032940E+1   2.032940E+1   -1.568000E+3   -1.568000E+3   8.999910E+1   -1.568000E+3   -1.568000E+3   -1.973917E-1   2.037039E-1   -4.186651E-4   -1.045128E-5   1.044471E-5   -4.186653E-4   4.187956E-4   -1.785700E+2   -8.857090E+1   
6.501984E+3   2.031021E+1   2.031021E+1   -1.579000E+3   -1.579000E+3   8.999910E+1   -1.578000E+3   -1.578000E+3   -1.959025E-1   2.064773E-1   -4.199957E-4   -1.348577E-5   1.347917E-5   -4.199959E-4   4.202121E-4   -1.781609E+2   -8.816180E+1   
6.528940E+3   2.030541E+1   2.030541E+1   -1.589000E+3   -1.589000E+3   8.999910E+1   -1.588000E+3   -1.588000E+3   -1.961025E-1   2.046134E-1   -4.195881E-4   -1.208565E-5   1.207906E-5   -4.195883E-4   4.197621E-4   -1.783501E+2   -8.835103E+1   
6.555888E+3   2.030941E+1   2.030941E+1   -1.598000E+3   -1.598000E+3   8.999910E+1   -1.597000E+3   -1.597000E+3   -1.956813E-1   2.047484E-1   -4.199401E-4   -1.251775E-5   1.251116E-5   -4.199403E-4   4.201266E-4   -1.782926E+2   -8.829351E+1   
6.582841E+3   2.032070E+1   2.032070E+1   -1.609000E+3   -1.609000E+3   8.999910E+1   -1.608000E+3   -1.608000E+3   -1.956585E-1   2.027980E-1   -4.193915E-4   -1.121652E-5   1.120993E-5   -4.193916E-4   4.195414E-4   -1.784680E+2   -8.846890E+1   
6.609847E+3   2.029510E+1   2.029510E+1   -1.619000E+3   -1.619000E+3   8.999910E+1   -1.618000E+3   -1.618000E+3   -1.930423E-1   2.014129E-1   -4.174000E-4   -1.210933E-5   1.210278E-5   -4.174002E-4   4.175757E-4   -1.783382E+2   -8.833914E+1   
6.636797E+3   2.030941E+1   2.030941E+1   -1.629000E+3   -1.629000E+3   8.999910E+1   -1.628000E+3   -1.628000E+3   -1.936118E-1   2.010189E-1   -4.181475E-4   -1.148619E-5   1.147962E-5   -4.181476E-4   4.183052E-4   -1.784265E+2   -8.842742E+1   
6.663712E+3   2.031741E+1   2.031741E+1   -1.638000E+3   -1.638000E+3   8.999910E+1   -1.638000E+3   -1.638000E+3   -1.928092E-1   1.991108E-1   -4.170434E-4   -1.075144E-5   1.074488E-5   -4.170436E-4   4.171820E-4   -1.785232E+2   -8.852413E+1   
6.691206E+3   2.032150E+1   2.032150E+1   -1.648000E+3   -1.648000E+3   8.999910E+1   -1.648000E+3   -1.648000E+3   -1.911152E-1   1.999511E-1   -4.170428E-4   -1.256874E-5   1.256219E-5   -4.170430E-4   4.172321E-4   -1.782738E+2   -8.827466E+1   
6.718141E+3   2.032559E+1   2.032559E+1   -1.658000E+3   -1.658000E+3   8.999910E+1   -1.657000E+3   -1.657000E+3   -1.905867E-1   1.968639E-1   -4.153320E-4   -1.080935E-5   1.080283E-5   -4.153321E-4   4.154726E-4   -1.785092E+2   -8.851007E+1   
6.745047E+3   2.032760E+1   2.032760E+1   -1.668000E+3   -1.668000E+3   8.999910E+1   -1.668000E+3   -1.668000E+3   -1.903694E-1   1.981108E-1   -4.166292E-4   -1.189175E-5   1.188520E-5   -4.166294E-4   4.167989E-4   -1.783651E+2   -8.836596E+1   
6.772513E+3   2.034481E+1   2.034481E+1   -1.678000E+3   -1.678000E+3   8.999910E+1   -1.678000E+3   -1.678000E+3   -1.900870E-1   1.980834E-1   -4.170345E-4   -1.211828E-5   1.211173E-5   -4.170347E-4   4.172105E-4   -1.783356E+2   -8.833646E+1   
6.799969E+3   2.035021E+1   2.035021E+1   -1.688000E+3   -1.688000E+3   8.999910E+1   -1.688000E+3   -1.688000E+3   -1.891866E-1   1.953581E-1   -4.153602E-4   -1.087670E-5   1.087017E-5   -4.153604E-4   4.155026E-4   -1.785000E+2   -8.850089E+1   
6.826969E+3   2.033260E+1   2.033260E+1   -1.698000E+3   -1.698000E+3   8.999910E+1   -1.698000E+3   -1.698000E+3   -1.890991E-1   1.972521E-1   -4.170829E-4   -1.231908E-5   1.231253E-5   -4.170831E-4   4.172648E-4   -1.783082E+2   -8.830909E+1   
6.853974E+3   2.035870E+1   2.035870E+1   -1.709000E+3   -1.709000E+3   8.999910E+1   -1.708000E+3   -1.708000E+3   -1.894047E-1   1.955305E-1   -4.168338E-4   -1.094559E-5   1.093904E-5   -4.168340E-4   4.169775E-4   -1.784958E+2   -8.849672E+1   
6.881690E+3   2.034301E+1   2.034301E+1   -1.718000E+3   -1.718000E+3   8.999910E+1   -1.718000E+3   -1.718000E+3   -1.861715E-1   1.964619E-1   -4.158621E-4   -1.389624E-5   1.388971E-5   -4.158623E-4   4.160942E-4   -1.780861E+2   -8.808704E+1   
6.908660E+3   2.034460E+1   2.034460E+1   -1.728000E+3   -1.728000E+3   8.999910E+1   -1.728000E+3   -1.728000E+3   -1.872236E-1   1.944064E-1   -4.159049E-4   -1.176939E-5   1.176286E-5   -4.159051E-4   4.160714E-4   -1.783791E+2   -8.837996E+1   
6.935607E+3   2.035909E+1   2.035909E+1   -1.738000E+3   -1.738000E+3   8.999910E+1   -1.738000E+3   -1.738000E+3   -1.885640E-1   1.975394E-1   -4.193462E-4   -1.309122E-5   1.308463E-5   -4.193464E-4   4.195505E-4   -1.782119E+2   -8.821281E+1   
6.962543E+3   2.034869E+1   2.034869E+1   -1.748000E+3   -1.748000E+3   8.999910E+1   -1.748000E+3   -1.748000E+3   -1.884583E-1   1.932945E-1   -4.172634E-4   -1.022894E-5   1.022239E-5   -4.172635E-4   4.173887E-4   -1.785957E+2   -8.859661E+1   
6.990786E+3   2.034240E+1   2.034240E+1   -1.758000E+3   -1.758000E+3   8.999910E+1   -1.757000E+3   -1.757000E+3   -1.834117E-1   1.909669E-1   -4.130064E-4   -1.214216E-5   1.213567E-5   -4.130066E-4   4.131849E-4   -1.783160E+2   -8.831692E+1   
7.017774E+3   2.033251E+1   2.033251E+1   -1.768000E+3   -1.768000E+3   8.999910E+1   -1.768000E+3   -1.768000E+3   -1.865789E-1   1.942434E-1   -4.178167E-4   -1.230096E-5   1.229440E-5   -4.178169E-4   4.179977E-4   -1.783136E+2   -8.831454E+1   
7.044802E+3   2.032400E+1   2.032400E+1   -1.778000E+3   -1.778000E+3   8.999910E+1   -1.778000E+3   -1.778000E+3   -1.857382E-1   1.945198E-1   -4.180371E-4   -1.312891E-5   1.312235E-5   -4.180373E-4   4.182432E-4   -1.782012E+2   -8.820205E+1   
7.073046E+3   2.032330E+1   2.032330E+1   -1.788000E+3   -1.788000E+3   8.999910E+1   -1.787000E+3   -1.787000E+3   -1.837433E-1   1.938559E-1   -4.168450E-4   -1.409241E-5   1.408587E-5   -4.168452E-4   4.170831E-4   -1.780637E+2   -8.806462E+1   
7.101337E+3   2.032629E+1   2.032629E+1   -1.798000E+3   -1.798000E+3   8.999910E+1   -1.797000E+3   -1.797000E+3   -1.845334E-1   1.911671E-1   -4.163216E-4   -1.170219E-5   1.169566E-5   -4.163218E-4   4.164861E-4   -1.783899E+2   -8.839082E+1   
7.128271E+3   2.032980E+1   2.032980E+1   -1.809000E+3   -1.809000E+3   8.999910E+1   -1.807000E+3   -1.807000E+3   -1.838740E-1   1.922106E-1   -4.171371E-4   -1.294374E-5   1.293719E-5   -4.171373E-4   4.173379E-4   -1.782227E+2   -8.822359E+1   
7.155220E+3   2.033019E+1   2.033019E+1   -1.818000E+3   -1.818000E+3   8.999910E+1   -1.817000E+3   -1.817000E+3   -1.831576E-1   1.906191E-1   -4.162862E-4   -1.237174E-5   1.236520E-5   -4.162864E-4   4.164700E-4   -1.782977E+2   -8.829861E+1   
7.182910E+3   2.030959E+1   2.030959E+1   -1.828000E+3   -1.828000E+3   8.999910E+1   -1.828000E+3   -1.828000E+3   -1.832731E-1   1.921275E-1   -4.179672E-4   -1.340687E-5   1.340031E-5   -4.179674E-4   4.181821E-4   -1.781628E+2   -8.816369E+1   
7.211195E+3   2.032131E+1   2.032131E+1   -1.838000E+3   -1.838000E+3   8.999910E+1   -1.837000E+3   -1.837000E+3   -1.857366E-1   1.932534E-1   -4.208568E-4   -1.253201E-5   1.252540E-5   -4.208570E-4   4.210434E-4   -1.782944E+2   -8.829529E+1   
7.238164E+3   2.031371E+1   2.031371E+1   -1.848000E+3   -1.848000E+3   8.999910E+1   -1.848000E+3   -1.848000E+3   -1.862873E-1   1.912350E-1   -4.206489E-4   -1.078460E-5   1.077799E-5   -4.206491E-4   4.207872E-4   -1.785314E+2   -8.853227E+1   
7.265095E+3   2.031671E+1   2.031671E+1   -1.858000E+3   -1.858000E+3   8.999910E+1   -1.857000E+3   -1.857000E+3   -1.834708E-1   1.925505E-1   -4.201316E-4   -1.371080E-5   1.370420E-5   -4.201318E-4   4.203553E-4   -1.781308E+2   -8.813174E+1   
7.293330E+3   2.033190E+1   2.033190E+1   -1.868000E+3   -1.868000E+3   8.999910E+1   -1.867000E+3   -1.867000E+3   -1.818373E-1   1.894524E-1   -4.177377E-4   -1.271636E-5   1.270979E-5   -4.177379E-4   4.179312E-4   -1.782564E+2   -8.825730E+1   
7.321608E+3   2.033981E+1   2.033981E+1   -1.878000E+3   -1.878000E+3   8.999910E+1   -1.877000E+3   -1.877000E+3   -1.807779E-1   1.879503E-1   -4.167131E-4   -1.244544E-5   1.243890E-5   -4.167133E-4   4.168989E-4   -1.782893E+2   -8.829023E+1   
7.348563E+3   2.034619E+1   2.034619E+1   -1.888000E+3   -1.888000E+3   8.999910E+1   -1.887000E+3   -1.887000E+3   -1.812697E-1   1.865270E-1   -4.167726E-4   -1.115246E-5   1.114591E-5   -4.167727E-4   4.169217E-4   -1.784672E+2   -8.846808E+1   
7.375509E+3   2.033941E+1   2.033941E+1   -1.898000E+3   -1.898000E+3   8.999910E+1   -1.897000E+3   -1.897000E+3   -1.814309E-1   1.861104E-1   -4.172335E-4   -1.079712E-5   1.079057E-5   -4.172336E-4   4.173732E-4   -1.785176E+2   -8.851854E+1   
7.403703E+3   2.034371E+1   2.034371E+1   -1.908000E+3   -1.908000E+3   8.999910E+1   -1.908000E+3   -1.908000E+3   -1.807227E-1   1.882114E-1   -4.187308E-4   -1.282115E-5   1.281457E-5   -4.187310E-4   4.189271E-4   -1.782462E+2   -8.824710E+1   
7.430693E+3   2.033181E+1   2.033181E+1   -1.918000E+3   -1.918000E+3   8.999910E+1   -1.917000E+3   -1.917000E+3   -1.797831E-1   1.874533E-1   -4.181849E-4   -1.298536E-5   1.297879E-5   -4.181851E-4   4.183864E-4   -1.782214E+2   -8.822234E+1   
7.457640E+3   2.032101E+1   2.032101E+1   -1.928000E+3   -1.928000E+3   8.999910E+1   -1.928000E+3   -1.928000E+3   -1.800024E-1   1.878592E-1   -4.192539E-4   -1.317296E-5   1.316637E-5   -4.192541E-4   4.194608E-4   -1.782004E+2   -8.820126E+1   
7.485305E+3   2.031631E+1   2.031631E+1   -1.938000E+3   -1.938000E+3   8.999910E+1   -1.937000E+3   -1.937000E+3   -1.799692E-1   1.870678E-1   -4.192924E-4   -1.268415E-5   1.267756E-5   -4.192926E-4   4.194842E-4   -1.782673E+2   -8.826816E+1   
7.513552E+3   2.032311E+1   2.032311E+1   -1.948000E+3   -1.948000E+3   8.999910E+1   -1.947000E+3   -1.947000E+3   -1.778780E-1   1.851443E-1   -4.173187E-4   -1.283358E-5   1.282703E-5   -4.173189E-4   4.175160E-4   -1.782386E+2   -8.823947E+1   
7.540596E+3   2.031771E+1   2.031771E+1   -1.958000E+3   -1.958000E+3   8.999910E+1   -1.957000E+3   -1.957000E+3   -1.785554E-1   1.839267E-1   -4.176292E-4   -1.155635E-5   1.154979E-5   -4.176294E-4   4.177890E-4   -1.784150E+2   -8.841585E+1   
7.567641E+3   2.030789E+1   2.030789E+1   -1.968000E+3   -1.968000E+3   8.999910E+1   -1.967000E+3   -1.967000E+3   -1.773491E-1   1.854795E-1   -4.183942E-4   -1.353598E-5   1.352940E-5   -4.183945E-4   4.186131E-4   -1.781470E+2   -8.814790E+1   
7.595843E+3   2.030740E+1   2.030740E+1   -1.978000E+3   -1.978000E+3   8.999910E+1   -1.977000E+3   -1.977000E+3   -1.762948E-1   1.849596E-1   -4.179800E-4   -1.395228E-5   1.394571E-5   -4.179803E-4   4.182128E-4   -1.780882E+2   -8.808906E+1   
7.624124E+3   2.029821E+1   2.029821E+1   -1.988000E+3   -1.988000E+3   8.999910E+1   -1.988000E+3   -1.988000E+3   -1.765995E-1   1.836381E-1   -4.180386E-4   -1.286583E-5   1.285926E-5   -4.180388E-4   4.182366E-4   -1.782372E+2   -8.823808E+1   
7.651110E+3   2.029949E+1   2.029949E+1   -1.998000E+3   -1.998000E+3   8.999910E+1   -1.997000E+3   -1.997000E+3   -1.762485E-1   1.825381E-1   -4.176743E-4   -1.238071E-5   1.237415E-5   -4.176745E-4   4.178577E-4   -1.783021E+2   -8.830303E+1   
7.692064E+3   2.030880E+1   2.030880E+1   -2.098000E+3   -2.098000E+3   8.999910E+1   -2.097000E+3   -2.097000E+3   -1.719976E-1   1.790140E-1   -4.187666E-4   -1.335112E-5   1.334454E-5   -4.187668E-4   4.189794E-4   -1.781739E+2   -8.817481E+1   
7.721005E+3   2.030840E+1   2.030840E+1   -2.198000E+3   -2.198000E+3   8.999910E+1   -2.198000E+3   -2.198000E+3   -1.681915E-1   1.749693E-1   -4.198953E-4   -1.365145E-5   1.364486E-5   -4.198955E-4   4.201171E-4   -1.781379E+2   -8.813878E+1   
7.749948E+3   2.029409E+1   2.029409E+1   -2.299000E+3   -2.299000E+3   8.999910E+1   -2.298000E+3   -2.298000E+3   -1.612730E-1   1.668853E-1   -4.163894E-4   -1.326807E-5   1.326153E-5   -4.163897E-4   4.166008E-4   -1.781749E+2   -8.817581E+1   
7.779692E+3   2.029571E+1   2.029571E+1   -2.398000E+3   -2.398000E+3   8.999910E+1   -2.398000E+3   -2.398000E+3   -1.584743E-1   1.576011E-1   -4.148918E-4   -9.178702E-6   9.172185E-6   -4.148919E-4   4.149933E-4   -1.787326E+2   -8.873355E+1   
7.808152E+3   2.029849E+1   2.029849E+1   -2.499000E+3   -2.499000E+3   8.999910E+1   -2.498000E+3   -2.498000E+3   -1.515458E-1   1.586645E-1   -4.170316E-4   -1.523548E-5   1.522893E-5   -4.170319E-4   4.173098E-4   -1.779077E+2   -8.790864E+1   
7.836556E+3   2.031841E+1   2.031841E+1   -2.599000E+3   -2.599000E+3   8.999910E+1   -2.598000E+3   -2.598000E+3   -1.473958E-1   1.536729E-1   -4.172845E-4   -1.510377E-5   1.509721E-5   -4.172847E-4   4.175578E-4   -1.779271E+2   -8.792796E+1   
7.866215E+3   2.031829E+1   2.031829E+1   -2.699000E+3   -2.699000E+3   8.999910E+1   -2.698000E+3   -2.698000E+3   -1.416348E-1   1.489485E-1   -4.166273E-4   -1.627903E-5   1.627249E-5   -4.166275E-4   4.169452E-4   -1.777624E+2   -8.776330E+1   
7.895132E+3   2.032549E+1   2.032549E+1   -2.799000E+3   -2.799000E+3   8.999910E+1   -2.798000E+3   -2.798000E+3   -1.382533E-1   1.411007E-1   -4.156282E-4   -1.360481E-5   1.359828E-5   -4.156284E-4   4.158508E-4   -1.781252E+2   -8.812610E+1   
7.923632E+3   2.034551E+1   2.034551E+1   -2.899000E+3   -2.899000E+3   8.999910E+1   -2.898000E+3   -2.898000E+3   -1.313238E-1   1.329808E-1   -4.120929E-4   -1.320377E-5   1.319730E-5   -4.120931E-4   4.123043E-4   -1.781648E+2   -8.816573E+1   
7.953264E+3   2.034460E+1   2.034460E+1   -2.999000E+3   -2.999000E+3   8.999910E+1   -2.998000E+3   -2.998000E+3   -1.265464E-1   1.327075E-1   -4.148425E-4   -1.682614E-5   1.681962E-5   -4.148428E-4   4.151836E-4   -1.776773E+2   -8.767824E+1   
7.982117E+3   2.032049E+1   2.032049E+1   -3.098000E+3   -3.098000E+3   8.999910E+1   -3.098000E+3   -3.098000E+3   -1.304490E-1   1.453945E-1   -4.313941E-4   -2.353372E-5   2.352695E-5   -4.313945E-4   4.320355E-4   -1.768775E+2   -8.687835E+1   
8.011057E+3   2.031979E+1   2.031979E+1   -3.198000E+3   -3.198000E+3   8.999910E+1   -3.197000E+3   -3.197000E+3   -1.276869E-1   1.383919E-1   -4.312696E-4   -2.101869E-5   2.101191E-5   -4.312700E-4   4.317815E-4   -1.772098E+2   -8.721070E+1   
8.040776E+3   2.033190E+1   2.033190E+1   -3.299000E+3   -3.299000E+3   8.999910E+1   -3.298000E+3   -3.298000E+3   -1.179704E-1   1.133871E-1   -4.155017E-4   -1.068384E-5   1.067731E-5   -4.155018E-4   4.156390E-4   -1.785271E+2   -8.852797E+1   
8.069720E+3   2.033129E+1   2.033129E+1   -3.398000E+3   -3.398000E+3   8.999910E+1   -3.398000E+3   -3.398000E+3   -1.122220E-1   1.165161E-1   -4.197055E-4   -1.737350E-5   1.736691E-5   -4.197058E-4   4.200649E-4   -1.776296E+2   -8.763052E+1   
8.098660E+3   2.033209E+1   2.033209E+1   -3.499000E+3   -3.499000E+3   8.999910E+1   -3.498000E+3   -3.498000E+3   -1.087633E-1   1.120044E-1   -4.207164E-4   -1.709906E-5   1.709245E-5   -4.207167E-4   4.210637E-4   -1.776726E+2   -8.767352E+1   
8.127857E+3   2.030999E+1   2.030999E+1   -3.598000E+3   -3.598000E+3   8.999910E+1   -3.597000E+3   -3.597000E+3   -1.040405E-1   1.077325E-1   -4.209706E-4   -1.786647E-5   1.785986E-5   -4.209709E-4   4.213495E-4   -1.775698E+2   -8.757066E+1   
8.157097E+3   2.030871E+1   2.030871E+1   -3.698000E+3   -3.698000E+3   8.999910E+1   -3.697000E+3   -3.697000E+3   -9.831320E-2   1.017463E-1   -4.195561E-4   -1.813094E-5   1.812435E-5   -4.195564E-4   4.199477E-4   -1.775255E+2   -8.752643E+1   
8.186331E+3   2.030029E+1   2.030029E+1   -3.798000E+3   -3.798000E+3   8.999910E+1   -3.797000E+3   -3.797000E+3   -9.403399E-2   9.803255E-2   -4.205124E-4   -1.898767E-5   1.898107E-5   -4.205127E-4   4.209408E-4   -1.774146E+2   -8.741554E+1   
8.215500E+3   2.029260E+1   2.029260E+1   -3.898000E+3   -3.898000E+3   8.999910E+1   -3.897000E+3   -3.897000E+3   -8.805756E-2   9.189370E-2   -4.188373E-4   -1.931786E-5   1.931128E-5   -4.188376E-4   4.192826E-4   -1.773592E+2   -8.736014E+1   
8.244681E+3   2.028149E+1   2.028149E+1   -3.998000E+3   -3.998000E+3   8.999910E+1   -3.997000E+3   -3.997000E+3   -8.550842E-2   9.029403E-2   -4.222546E-4   -2.045959E-5   2.045295E-5   -4.222550E-4   4.227500E-4   -1.772260E+2   -8.722691E+1   
8.274349E+3   2.028149E+1   2.028149E+1   -4.098000E+3   -4.098000E+3   8.999910E+1   -4.097000E+3   -4.097000E+3   -8.022123E-2   8.430761E-2   -4.211338E-4   -2.041819E-5   2.041157E-5   -4.211341E-4   4.216285E-4   -1.772243E+2   -8.722515E+1   
8.303601E+3   2.027950E+1   2.027950E+1   -4.198000E+3   -4.198000E+3   8.999910E+1   -4.198000E+3   -4.198000E+3   -7.535514E-2   7.933883E-2   -4.209839E-4   -2.080493E-5   2.079831E-5   -4.209842E-4   4.214977E-4   -1.771708E+2   -8.717166E+1   
8.332494E+3   2.029031E+1   2.029031E+1   -4.298000E+3   -4.298000E+3   8.999910E+1   -4.298000E+3   -4.298000E+3   -6.898907E-2   7.160036E-2   -4.180603E-4   -2.028079E-5   2.027422E-5   -4.180606E-4   4.185520E-4   -1.772227E+2   -8.722357E+1   
8.360948E+3   2.029351E+1   2.029351E+1   -4.399000E+3   -4.399000E+3   8.999910E+1   -4.398000E+3   -4.398000E+3   -6.520593E-2   7.076549E-2   -4.211266E-4   -2.281758E-5   2.281097E-5   -4.211269E-4   4.217443E-4   -1.768986E+2   -8.689952E+1   
8.390193E+3   2.030410E+1   2.030410E+1   -4.499000E+3   -4.499000E+3   8.999910E+1   -4.498000E+3   -4.498000E+3   -5.913905E-2   6.557188E-2   -4.199752E-4   -2.387536E-5   2.386876E-5   -4.199756E-4   4.206533E-4   -1.767463E+2   -8.674717E+1   
8.418598E+3   2.029379E+1   2.029379E+1   -4.599000E+3   -4.599000E+3   8.999910E+1   -4.598000E+3   -4.598000E+3   -5.541896E-2   5.910188E-2   -4.196015E-4   -2.240529E-5   2.239870E-5   -4.196019E-4   4.201993E-4   -1.769435E+2   -8.694440E+1   
8.446497E+3   2.031481E+1   2.031481E+1   -4.699000E+3   -4.699000E+3   8.999910E+1   -4.699000E+3   -4.699000E+3   -5.068117E-2   5.209192E-2   -4.182760E-4   -2.126738E-5   2.126081E-5   -4.182763E-4   4.188163E-4   -1.770893E+2   -8.709018E+1   
8.475740E+3   2.031201E+1   2.031201E+1   -4.799000E+3   -4.799000E+3   8.999910E+1   -4.798000E+3   -4.798000E+3   -4.193534E-2   4.548296E-2   -4.144009E-4   -2.318574E-5   2.317923E-5   -4.144013E-4   4.150490E-4   -1.767976E+2   -8.679854E+1   
8.503724E+3   2.029641E+1   2.029641E+1   -4.899000E+3   -4.899000E+3   8.999910E+1   -4.898000E+3   -4.898000E+3   -3.739621E-2   4.483397E-2   -4.170774E-4   -2.637841E-5   2.637186E-5   -4.170779E-4   4.179108E-4   -1.763811E+2   -8.638200E+1   
8.531712E+3   2.030761E+1   2.030761E+1   -4.999000E+3   -4.999000E+3   8.999910E+1   -4.998000E+3   -4.998000E+3   -3.060932E-2   4.212242E-2   -4.169792E-4   -2.968192E-5   2.967537E-5   -4.169797E-4   4.180343E-4   -1.759284E+2   -8.592927E+1   
8.560641E+3   2.029312E+1   2.029312E+1   -5.099000E+3   -5.099000E+3   8.999910E+1   -5.099000E+3   -5.099000E+3   -2.888593E-2   3.330684E-2   -4.165499E-4   -2.518021E-5   2.517367E-5   -4.165503E-4   4.173103E-4   -1.765407E+2   -8.654161E+1   
8.589095E+3   2.030959E+1   2.030959E+1   -5.199000E+3   -5.199000E+3   8.999910E+1   -5.198000E+3   -5.198000E+3   -2.466977E-2   2.817841E-2   -4.166130E-4   -2.499327E-5   2.498673E-5   -4.166134E-4   4.173620E-4   -1.765669E+2   -8.656775E+1   
8.617062E+3   2.031161E+1   2.031161E+1   -5.299000E+3   -5.299000E+3   8.999910E+1   -5.298000E+3   -5.298000E+3   -1.844200E-2   2.241163E-2   -4.150001E-4   -2.575971E-5   2.575320E-5   -4.150005E-4   4.157988E-4   -1.764481E+2   -8.644902E+1   
8.646808E+3   2.030059E+1   2.030059E+1   -5.399000E+3   -5.399000E+3   8.999910E+1   -5.398000E+3   -5.398000E+3   -1.536148E-2   2.058467E-2   -4.179223E-4   -2.711072E-5   2.710415E-5   -4.179227E-4   4.188007E-4   -1.762884E+2   -8.628931E+1   
8.675267E+3   2.029821E+1   2.029821E+1   -5.499000E+3   -5.499000E+3   8.999910E+1   -5.498000E+3   -5.498000E+3   -1.095429E-2   1.372464E-2   -4.168490E-4   -2.584364E-5   2.583709E-5   -4.168494E-4   4.176493E-4   -1.764523E+2   -8.645324E+1   
8.703193E+3   2.032961E+1   2.032961E+1   -5.599000E+3   -5.599000E+3   8.999910E+1   -5.598000E+3   -5.598000E+3   -1.273951E-3   4.834381E-3   -4.110016E-4   -2.681173E-5   2.680527E-5   -4.110020E-4   4.118752E-4   -1.762676E+2   -8.626849E+1   
8.732449E+3   2.031719E+1   2.031719E+1   -5.699000E+3   -5.699000E+3   8.999910E+1   -5.698000E+3   -5.698000E+3   2.532363E-3   7.353951E-3   -4.161252E-4   -3.172372E-5   3.171719E-5   -4.161257E-4   4.173327E-4   -1.756404E+2   -8.564133E+1   
8.760897E+3   2.031030E+1   2.031030E+1   -5.799000E+3   -5.799000E+3   8.999910E+1   -5.798000E+3   -5.798000E+3   4.284395E-3   -5.145476E-3   -4.133394E-4   -2.464618E-5   2.463969E-5   -4.133397E-4   4.140735E-4   -1.765877E+2   -8.658857E+1   
8.789354E+3   2.029931E+1   2.029931E+1   -5.899000E+3   -5.899000E+3   8.999910E+1   -5.898000E+3   -5.898000E+3   1.166546E-2   -1.253081E-2   -4.099565E-4   -2.507547E-5   2.506903E-5   -4.099569E-4   4.107227E-4   -1.764998E+2   -8.650070E+1   
8.819048E+3   2.030151E+1   2.030151E+1   -5.999000E+3   -5.999000E+3   8.999910E+1   -5.998000E+3   -5.998000E+3   1.739446E-2   -1.443611E-2   -4.110626E-4   -2.821113E-5   2.820468E-5   -4.110630E-4   4.120295E-4   -1.760740E+2   -8.607486E+1   
8.858345E+3   2.030691E+1   2.030691E+1   -5.899000E+3   -5.899000E+3   8.999910E+1   -5.898000E+3   -5.898000E+3   1.067153E-2   -7.758592E-3   -4.135688E-4   -2.774123E-5   2.773473E-5   -4.135692E-4   4.144981E-4   -1.761625E+2   -8.616338E+1   
8.885522E+3   2.029180E+1   2.029180E+1   -5.799000E+3   -5.799000E+3   8.999910E+1   -5.798000E+3   -5.798000E+3   5.962992E-3   -4.302067E-3   -4.127401E-4   -2.640537E-5   2.639888E-5   -4.127405E-4   4.135839E-4   -1.763394E+2   -8.634035E+1   
8.912471E+3   2.029669E+1   2.029669E+1   -5.699000E+3   -5.699000E+3   8.999910E+1   -5.698000E+3   -5.698000E+3   2.299270E-3   1.777622E-3   -4.128350E-4   -2.764010E-5   2.763361E-5   -4.128355E-4   4.137593E-4   -1.761697E+2   -8.617055E+1   
8.939377E+3   2.029449E+1   2.029449E+1   -5.599000E+3   -5.599000E+3   8.999910E+1   -5.598000E+3   -5.598000E+3   -3.653665E-3   6.392006E-3   -4.135524E-4   -2.625411E-5   2.624761E-5   -4.135528E-4   4.143849E-4   -1.763675E+2   -8.636839E+1   
8.966334E+3   2.030471E+1   2.030471E+1   -5.498000E+3   -5.498000E+3   8.999910E+1   -5.498000E+3   -5.498000E+3   -9.808921E-3   1.059566E-2   -4.141511E-4   -2.443873E-5   2.443222E-5   -4.141514E-4   4.148715E-4   -1.766229E+2   -8.662384E+1   
8.993249E+3   2.029559E+1   2.029559E+1   -5.399000E+3   -5.399000E+3   8.999910E+1   -5.398000E+3   -5.398000E+3   -1.473654E-2   1.669973E-2   -4.151046E-4   -2.481264E-5   2.480612E-5   -4.151050E-4   4.158455E-4   -1.765792E+2   -8.658015E+1   
9.020480E+3   2.030169E+1   2.030169E+1   -5.299000E+3   -5.299000E+3   8.999910E+1   -5.299000E+3   -5.299000E+3   -1.829453E-2   2.201675E-2   -4.147187E-4   -2.558941E-5   2.558289E-5   -4.147191E-4   4.155075E-4   -1.764692E+2   -8.647005E+1   
9.047664E+3   2.031451E+1   2.031451E+1   -5.199000E+3   -5.199000E+3   8.999910E+1   -5.198000E+3   -5.198000E+3   -2.432547E-2   2.528801E-2   -4.145972E-4   -2.319968E-5   2.319317E-5   -4.145976E-4   4.152458E-4   -1.767972E+2   -8.679813E+1   
9.074603E+3   2.031979E+1   2.031979E+1   -5.099000E+3   -5.099000E+3   8.999910E+1   -5.098000E+3   -5.098000E+3   -2.829266E-2   3.128211E-2   -4.148417E-4   -2.416342E-5   2.415690E-5   -4.148421E-4   4.155449E-4   -1.766664E+2   -8.666734E+1   
9.101788E+3   2.032198E+1   2.032198E+1   -4.999000E+3   -4.999000E+3   8.999910E+1   -4.998000E+3   -4.998000E+3   -3.384096E-2   3.884600E-2   -4.171116E-4   -2.513283E-5   2.512628E-5   -4.171120E-4   4.178681E-4   -1.765518E+2   -8.655274E+1   
9.128987E+3   2.032198E+1   2.032198E+1   -4.899000E+3   -4.899000E+3   8.999910E+1   -4.898000E+3   -4.898000E+3   -3.774967E-2   4.162302E-2   -4.153293E-4   -2.387469E-5   2.386817E-5   -4.153296E-4   4.160149E-4   -1.767100E+2   -8.671094E+1   
9.155950E+3   2.032739E+1   2.032739E+1   -4.799000E+3   -4.799000E+3   8.999910E+1   -4.798000E+3   -4.798000E+3   -4.286650E-2   4.711066E-2   -4.160282E-4   -2.368364E-5   2.367711E-5   -4.160286E-4   4.167018E-4   -1.767418E+2   -8.674268E+1   
9.183245E+3   2.032839E+1   2.032839E+1   -4.699000E+3   -4.699000E+3   8.999910E+1   -4.698000E+3   -4.698000E+3   -4.833984E-2   5.206296E-2   -4.166343E-4   -2.286845E-5   2.286190E-5   -4.166346E-4   4.172614E-4   -1.768583E+2   -8.685917E+1   
9.210486E+3   2.033331E+1   2.033331E+1   -4.599000E+3   -4.599000E+3   8.999910E+1   -4.598000E+3   -4.598000E+3   -5.450486E-2   5.717434E-2   -4.178003E-4   -2.168467E-5   2.167810E-5   -4.178007E-4   4.183627E-4   -1.770289E+2   -8.702980E+1   
9.237423E+3   2.034069E+1   2.034069E+1   -4.499000E+3   -4.499000E+3   8.999910E+1   -4.498000E+3   -4.498000E+3   -5.860065E-2   6.220038E-2   -4.175326E-4   -2.187825E-5   2.187169E-5   -4.175329E-4   4.181054E-4   -1.770005E+2   -8.700141E+1   
9.264352E+3   2.032180E+1   2.032180E+1   -4.399000E+3   -4.399000E+3   8.999910E+1   -4.398000E+3   -4.398000E+3   -6.261995E-2   6.880960E-2   -4.181920E-4   -2.323839E-5   2.323183E-5   -4.181924E-4   4.188372E-4   -1.768194E+2   -8.682032E+1   
9.291299E+3   2.033111E+1   2.033111E+1   -4.299000E+3   -4.299000E+3   8.999910E+1   -4.298000E+3   -4.298000E+3   -7.007501E-2   7.526836E-2   -4.210517E-4   -2.210606E-5   2.209945E-5   -4.210520E-4   4.216316E-4   -1.769946E+2   -8.699552E+1   
9.318220E+3   2.034670E+1   2.034670E+1   -4.198000E+3   -4.198000E+3   8.999910E+1   -4.198000E+3   -4.198000E+3   -7.512786E-2   7.618882E-2   -4.188857E-4   -1.874747E-5   1.874089E-5   -4.188860E-4   4.193051E-4   -1.774374E+2   -8.743831E+1   
9.345130E+3   2.034261E+1   2.034261E+1   -4.098000E+3   -4.098000E+3   8.999910E+1   -4.097000E+3   -4.097000E+3   -7.706303E-2   8.246294E-2   -4.178860E-4   -2.131471E-5   2.130815E-5   -4.178863E-4   4.184292E-4   -1.770801E+2   -8.708100E+1   
9.372065E+3   2.035549E+1   2.035549E+1   -3.998000E+3   -3.998000E+3   8.999910E+1   -3.998000E+3   -3.998000E+3   -8.753531E-2   8.800393E-2   -4.222535E-4   -1.744599E-5   1.743936E-5   -4.222537E-4   4.226137E-4   -1.776341E+2   -8.763499E+1   
9.399240E+3   2.036639E+1   2.036639E+1   -3.898000E+3   -3.898000E+3   8.999910E+1   -3.898000E+3   -3.898000E+3   -8.744385E-2   9.575828E-2   -4.208768E-4   -2.246701E-5   2.246039E-5   -4.208771E-4   4.214760E-4   -1.769444E+2   -8.694527E+1   
9.426455E+3   2.036480E+1   2.036480E+1   -3.798000E+3   -3.798000E+3   8.999910E+1   -3.797000E+3   -3.797000E+3   -9.216218E-2   1.017938E-1   -4.215872E-4   -2.293312E-5   2.292650E-5   -4.215875E-4   4.222105E-4   -1.768863E+2   -8.688724E+1   
9.453427E+3   2.035131E+1   2.035131E+1   -3.698000E+3   -3.698000E+3   8.999910E+1   -3.698000E+3   -3.698000E+3   -9.947294E-2   1.020528E-1   -4.205807E-4   -1.754585E-5   1.753924E-5   -4.205809E-4   4.209465E-4   -1.776111E+2   -8.761201E+1   
9.480599E+3   2.035269E+1   2.035269E+1   -3.598000E+3   -3.598000E+3   8.999910E+1   -3.598000E+3   -3.598000E+3   -1.059753E-1   1.106558E-1   -4.241294E-4   -1.858332E-5   1.857665E-5   -4.241297E-4   4.245363E-4   -1.774912E+2   -8.749208E+1   
9.507789E+3   2.035079E+1   2.035079E+1   -3.499000E+3   -3.499000E+3   8.999910E+1   -3.498000E+3   -3.498000E+3   -1.099510E-1   1.156788E-1   -4.237796E-4   -1.885814E-5   1.885148E-5   -4.237799E-4   4.241990E-4   -1.774520E+2   -8.745293E+1   
9.534977E+3   2.034820E+1   2.034820E+1   -3.399000E+3   -3.399000E+3   8.999910E+1   -3.398000E+3   -3.398000E+3   -1.133362E-1   1.197319E-1   -4.224363E-4   -1.886107E-5   1.885444E-5   -4.224366E-4   4.228572E-4   -1.774435E+2   -8.744444E+1   
9.561971E+3   2.034219E+1   2.034219E+1   -3.299000E+3   -3.299000E+3   8.999910E+1   -3.298000E+3   -3.298000E+3   -1.181855E-1   1.242438E-1   -4.223538E-4   -1.816973E-5   1.816309E-5   -4.223541E-4   4.227445E-4   -1.775366E+2   -8.753755E+1   
9.589135E+3   2.033569E+1   2.033569E+1   -3.198000E+3   -3.198000E+3   8.999910E+1   -3.198000E+3   -3.198000E+3   -1.235738E-1   1.292177E-1   -4.229165E-4   -1.742881E-5   1.742216E-5   -4.229167E-4   4.232755E-4   -1.776401E+2   -8.764102E+1   
9.616333E+3   2.034789E+1   2.034789E+1   -3.099000E+3   -3.099000E+3   8.999910E+1   -3.098000E+3   -3.098000E+3   -1.284301E-1   1.353736E-1   -4.238544E-4   -1.788868E-5   1.788202E-5   -4.238547E-4   4.242317E-4   -1.775833E+2   -8.758418E+1   
9.643517E+3   2.034539E+1   2.034539E+1   -2.999000E+3   -2.999000E+3   8.999910E+1   -2.998000E+3   -2.998000E+3   -1.331935E-1   1.388526E-1   -4.230763E-4   -1.653057E-5   1.652392E-5   -4.230765E-4   4.233991E-4   -1.777625E+2   -8.776336E+1   
9.670725E+3   2.033792E+1   2.033792E+1   -2.899000E+3   -2.899000E+3   8.999910E+1   -2.899000E+3   -2.899000E+3   -1.385461E-1   1.458071E-1   -4.249001E-4   -1.721225E-5   1.720557E-5   -4.249003E-4   4.252485E-4   -1.776803E+2   -8.768118E+1   
9.697973E+3   2.035760E+1   2.035760E+1   -2.799000E+3   -2.799000E+3   8.999910E+1   -2.798000E+3   -2.798000E+3   -1.469403E-1   1.517076E-1   -4.279805E-4   -1.503001E-5   1.502329E-5   -4.279807E-4   4.282443E-4   -1.779887E+2   -8.798959E+1   
9.724904E+3   2.035940E+1   2.035940E+1   -2.699000E+3   -2.699000E+3   8.999910E+1   -2.698000E+3   -2.698000E+3   -1.496899E-1   1.575746E-1   -4.273338E-4   -1.675014E-5   1.674343E-5   -4.273341E-4   4.276620E-4   -1.777553E+2   -8.775624E+1   
9.752045E+3   2.037640E+1   2.037640E+1   -2.599000E+3   -2.599000E+3   8.999910E+1   -2.598000E+3   -2.598000E+3   -1.517115E-1   1.575919E-1   -4.225867E-4   -1.486203E-5   1.485539E-5   -4.225869E-4   4.228480E-4   -1.779858E+2   -8.798668E+1   
9.779527E+3   2.037649E+1   2.037649E+1   -2.499000E+3   -2.499000E+3   8.999910E+1   -2.499000E+3   -2.499000E+3   -1.603138E-1   1.696989E-1   -4.297633E-4   -1.691005E-5   1.690329E-5   -4.297636E-4   4.300959E-4   -1.777467E+2   -8.774763E+1   
9.806504E+3   2.037600E+1   2.037600E+1   -2.399000E+3   -2.399000E+3   8.999910E+1   -2.398000E+3   -2.398000E+3   -1.626765E-1   1.698717E-1   -4.252788E-4   -1.488938E-5   1.488270E-5   -4.252790E-4   4.255393E-4   -1.779948E+2   -8.799574E+1   
9.833656E+3   2.038659E+1   2.038659E+1   -2.299000E+3   -2.299000E+3   8.999910E+1   -2.298000E+3   -2.298000E+3   -1.686702E-1   1.788482E-1   -4.287188E-4   -1.654287E-5   1.653613E-5   -4.287191E-4   4.290379E-4   -1.777902E+2   -8.779114E+1   
9.860897E+3   2.039059E+1   2.039059E+1   -2.199000E+3   -2.199000E+3   8.999910E+1   -2.198000E+3   -2.198000E+3   -1.730073E-1   1.816366E-1   -4.272294E-4   -1.499505E-5   1.498834E-5   -4.272296E-4   4.274925E-4   -1.779898E+2   -8.799074E+1   
9.888088E+3   2.040389E+1   2.040389E+1   -2.098000E+3   -2.098000E+3   8.999910E+1   -2.098000E+3   -2.098000E+3   -1.772711E-1   1.845589E-1   -4.257738E-4   -1.359250E-5   1.358581E-5   -4.257740E-4   4.259907E-4   -1.781715E+2   -8.817240E+1   
9.915240E+3   2.041161E+1   2.041161E+1   -1.998000E+3   -1.998000E+3   8.999910E+1   -1.998000E+3   -1.998000E+3   -1.812922E-1   1.909446E-1   -4.262964E-4   -1.479416E-5   1.478747E-5   -4.262966E-4   4.265530E-4   -1.780124E+2   -8.801331E+1   
9.954063E+3   2.040539E+1   2.040539E+1   -1.948000E+3   -1.948000E+3   8.999910E+1   -1.948000E+3   -1.948000E+3   -1.859874E-1   1.945027E-1   -4.285752E-4   -1.378696E-5   1.378022E-5   -4.285754E-4   4.287969E-4   -1.781575E+2   -8.815837E+1   
9.981191E+3   2.041421E+1   2.041421E+1   -1.898000E+3   -1.898000E+3   8.999910E+1   -1.897000E+3   -1.897000E+3   -1.877803E-1   1.958035E-1   -4.274610E-4   -1.320341E-5   1.319669E-5   -4.274612E-4   4.276648E-4   -1.782308E+2   -8.823171E+1   
1.000820E+4   2.042730E+1   2.042730E+1   -1.849000E+3   -1.849000E+3   8.999910E+1   -1.848000E+3   -1.848000E+3   -1.911324E-1   2.005831E-1   -4.296592E-4   -1.399327E-5   1.398652E-5   -4.296594E-4   4.298870E-4   -1.781346E+2   -8.813553E+1   
1.003516E+4   2.041329E+1   2.041329E+1   -1.798000E+3   -1.798000E+3   8.999910E+1   -1.798000E+3   -1.798000E+3   -1.937739E-1   2.030555E-1   -4.298964E-4   -1.364912E-5   1.364237E-5   -4.298966E-4   4.301130E-4   -1.781815E+2   -8.818238E+1   
1.006233E+4   2.042681E+1   2.042681E+1   -1.749000E+3   -1.749000E+3   8.999910E+1   -1.748000E+3   -1.748000E+3   -1.950717E-1   2.050559E-1   -4.289451E-4   -1.390642E-5   1.389968E-5   -4.289453E-4   4.291705E-4   -1.781431E+2   -8.814402E+1   
1.008953E+4   2.041812E+1   2.041812E+1   -1.699000E+3   -1.699000E+3   8.999910E+1   -1.698000E+3   -1.698000E+3   -1.994250E-1   2.068743E-1   -4.299208E-4   -1.191328E-5   1.190653E-5   -4.299209E-4   4.300858E-4   -1.784127E+2   -8.841362E+1   
1.011648E+4   2.042410E+1   2.042410E+1   -1.649000E+3   -1.649000E+3   8.999910E+1   -1.648000E+3   -1.648000E+3   -2.005781E-1   2.088104E-1   -4.288331E-4   -1.222596E-5   1.221923E-5   -4.288333E-4   4.290073E-4   -1.783669E+2   -8.836785E+1   
1.014342E+4   2.043279E+1   2.043279E+1   -1.598000E+3   -1.598000E+3   8.999910E+1   -1.598000E+3   -1.598000E+3   -2.021674E-1   2.115277E-1   -4.285193E-4   -1.278497E-5   1.277824E-5   -4.285195E-4   4.287100E-4   -1.782911E+2   -8.829197E+1   
1.017036E+4   2.043719E+1   2.043719E+1   -1.548000E+3   -1.548000E+3   8.999910E+1   -1.548000E+3   -1.548000E+3   -2.049057E-1   2.121499E-1   -4.276779E-4   -1.107238E-5   1.106566E-5   -4.276780E-4   4.278212E-4   -1.785170E+2   -8.851787E+1   
1.019725E+4   2.043691E+1   2.043691E+1   -1.499000E+3   -1.499000E+3   8.999910E+1   -1.498000E+3   -1.498000E+3   -2.053837E-1   2.164888E-1   -4.276244E-4   -1.354376E-5   1.353704E-5   -4.276247E-4   4.278389E-4   -1.781859E+2   -8.818683E+1   
1.022449E+4   2.043060E+1   2.043060E+1   -1.449000E+3   -1.449000E+3   8.999910E+1   -1.448000E+3   -1.448000E+3   -2.074005E-1   2.177216E-1   -4.266787E-4   -1.276181E-5   1.275511E-5   -4.266789E-4   4.268695E-4   -1.782868E+2   -8.828771E+1   
1.025166E+4   2.041509E+1   2.041509E+1   -1.399000E+3   -1.399000E+3   8.999910E+1   -1.398000E+3   -1.398000E+3   -2.104695E-1   2.190096E-1   -4.264693E-4   -1.128778E-5   1.128108E-5   -4.264695E-4   4.266187E-4   -1.784839E+2   -8.848475E+1   
1.027865E+4   2.043081E+1   2.043081E+1   -1.349000E+3   -1.349000E+3   8.999910E+1   -1.349000E+3   -1.349000E+3   -2.119634E-1   2.209947E-1   -4.257006E-4   -1.140307E-5   1.139638E-5   -4.257008E-4   4.258533E-4   -1.784656E+2   -8.846651E+1   
1.030558E+4   2.042449E+1   2.042449E+1   -1.299000E+3   -1.299000E+3   8.999910E+1   -1.299000E+3   -1.299000E+3   -2.164312E-1   2.269759E-1   -4.293249E-4   -1.225801E-5   1.225126E-5   -4.293251E-4   4.294999E-4   -1.783645E+2   -8.836545E+1   
1.033256E+4   2.042639E+1   2.042639E+1   -1.249000E+3   -1.249000E+3   8.999910E+1   -1.249000E+3   -1.249000E+3   -2.176430E-1   2.287374E-1   -4.281686E-4   -1.240706E-5   1.240034E-5   -4.281688E-4   4.283483E-4   -1.783402E+2   -8.834110E+1   
1.035944E+4   2.042120E+1   2.042120E+1   -1.199000E+3   -1.199000E+3   8.999910E+1   -1.199000E+3   -1.199000E+3   -2.209606E-1   2.308648E-1   -4.286439E-4   -1.135068E-5   1.134395E-5   -4.286440E-4   4.287941E-4   -1.784831E+2   -8.848404E+1   
1.038662E+4   2.042730E+1   2.042730E+1   -1.149000E+3   -1.149000E+3   8.999910E+1   -1.149000E+3   -1.149000E+3   -2.229908E-1   2.331900E-1   -4.283821E-4   -1.132762E-5   1.132090E-5   -4.283822E-4   4.285318E-4   -1.784853E+2   -8.848619E+1   
1.041357E+4   2.042571E+1   2.042571E+1   -1.099000E+3   -1.099000E+3   8.999910E+1   -1.099000E+3   -1.099000E+3   -2.257148E-1   2.376852E-1   -4.299243E-4   -1.234880E-5   1.234205E-5   -4.299245E-4   4.301016E-4   -1.783547E+2   -8.835563E+1   
1.044050E+4   2.041589E+1   2.041589E+1   -1.050000E+3   -1.050000E+3   8.999910E+1   -1.049000E+3   -1.049000E+3   -2.280150E-1   2.386773E-1   -4.290190E-4   -1.120073E-5   1.119399E-5   -4.290192E-4   4.291652E-4   -1.785045E+2   -8.850538E+1   
1.046765E+4   2.042629E+1   2.042629E+1   -9.990000E+2   -9.990000E+2   8.999910E+1   -9.990000E+2   -9.990000E+2   -2.304913E-1   2.413139E-1   -4.292474E-4   -1.108682E-5   1.108008E-5   -4.292475E-4   4.293905E-4   -1.785205E+2   -8.852136E+1   
1.049449E+4   2.042990E+1   2.042990E+1   -9.500000E+2   -9.500000E+2   8.999910E+1   -9.490000E+2   -9.490000E+2   -2.317893E-1   2.418336E-1   -4.273813E-4   -1.030270E-5   1.029599E-5   -4.273815E-4   4.275055E-4   -1.786191E+2   -8.861996E+1   
1.052126E+4   2.041839E+1   2.041839E+1   -9.000000E+2   -9.000000E+2   8.999910E+1   -8.990000E+2   -8.990000E+2   -2.117294E-1   2.196162E-1   -3.972101E-4   -8.364231E-6   8.357992E-6   -3.972103E-4   3.972982E-4   -1.787937E+2   -8.879458E+1   
1.054806E+4   2.042150E+1   2.042150E+1   -8.500000E+2   -8.500000E+2   8.999910E+1   -8.490000E+2   -8.490000E+2   -1.428125E-1   1.434335E-1   -3.010831E-4   -2.411571E-6   2.406842E-6   -3.010831E-4   3.010927E-4   -1.795411E+2   -8.954199E+1   
1.057486E+4   2.042349E+1   2.042349E+1   -7.990000E+2   -7.990000E+2   8.999910E+1   -7.990000E+2   -7.990000E+2   -1.177065E-1   1.178065E-1   -2.654370E-4   -1.580459E-6   1.576290E-6   -2.654371E-4   2.654417E-4   -1.796589E+2   -8.965975E+1   
1.060170E+4   2.043429E+1   2.043429E+1   -7.500000E+2   -7.500000E+2   8.999910E+1   -7.490000E+2   -7.490000E+2   -1.021288E-1   9.911031E-2   -2.404334E-4   9.951081E-7   -9.988849E-7   -2.404333E-4   2.404354E-4   1.797629E+2   2.697620E+2   
1.062845E+4   2.042840E+1   2.042840E+1   -7.000000E+2   -7.000000E+2   8.999910E+1   -6.990000E+2   -6.990000E+2   -8.850386E-2   8.504134E-2   -2.195923E-4   1.672969E-6   -1.676418E-6   -2.195922E-4   2.195986E-4   1.795635E+2   2.695626E+2   
1.065530E+4   2.042590E+1   2.042590E+1   -6.500000E+2   -6.500000E+2   8.999910E+1   -6.490000E+2   -6.490000E+2   -7.572293E-2   7.074809E-2   -1.991759E-4   3.094845E-6   -3.097974E-6   -1.991759E-4   1.992000E-4   1.791098E+2   2.691089E+2   
1.068207E+4   2.043191E+1   2.043191E+1   -5.990000E+2   -5.990000E+2   8.999910E+1   -5.990000E+2   -5.990000E+2   -6.511484E-2   6.042396E-2   -1.826625E-4   3.234689E-6   -3.237558E-6   -1.826624E-4   1.826911E-4   1.789855E+2   2.689846E+2   
1.070895E+4   2.044970E+1   2.044970E+1   -5.500000E+2   -5.500000E+2   8.999910E+1   -5.490000E+2   -5.490000E+2   -5.444212E-2   5.244264E-2   -1.675535E-4   1.681990E-6   -1.684622E-6   -1.675535E-4   1.675620E-4   1.794249E+2   2.694240E+2   
1.073567E+4   2.045281E+1   2.045281E+1   -4.990000E+2   -4.990000E+2   8.999910E+1   -4.990000E+2   -4.990000E+2   -4.562861E-2   4.269161E-2   -1.525920E-4   2.665382E-6   -2.667779E-6   -1.525920E-4   1.526153E-4   1.789993E+2   2.689984E+2   
1.076253E+4   2.044930E+1   2.044930E+1   -4.490000E+2   -4.490000E+2   8.999910E+1   -4.490000E+2   -4.490000E+2   -3.777218E-2   3.362403E-2   -1.386916E-4   3.832963E-6   -3.835141E-6   -1.386915E-4   1.387445E-4   1.784169E+2   2.684160E+2   
1.078929E+4   2.046240E+1   2.046240E+1   -3.990000E+2   -3.990000E+2   8.999910E+1   -3.980000E+2   -3.980000E+2   -2.997799E-2   2.764242E-2   -1.266785E-4   2.878431E-6   -2.880421E-6   -1.266785E-4   1.267112E-4   1.786983E+2   2.686974E+2   
1.081610E+4   2.042669E+1   2.042669E+1   -3.490000E+2   -3.490000E+2   8.999910E+1   -3.490000E+2   -3.490000E+2   -2.051304E-2   1.889449E-2   -1.119631E-4   2.698884E-6   -2.700643E-6   -1.119630E-4   1.119956E-4   1.786191E+2   2.686182E+2   
1.084288E+4   2.043109E+1   2.043109E+1   -2.990000E+2   -2.990000E+2   8.999910E+1   -2.990000E+2   -2.990000E+2   -1.360671E-2   1.287056E-2   -1.005775E-4   2.385913E-6   -2.387493E-6   -1.005775E-4   1.006058E-4   1.786411E+2   2.686402E+2   
1.086971E+4   2.043649E+1   2.043649E+1   -2.490000E+2   -2.490000E+2   8.999910E+1   -2.490000E+2   -2.490000E+2   -6.592503E-3   5.730198E-3   -8.843009E-5   2.783163E-6   -2.784552E-6   -8.843005E-5   8.847388E-5   1.781973E+2   2.681964E+2   
1.089645E+4   2.043191E+1   2.043191E+1   -1.990000E+2   -1.990000E+2   8.999910E+1   -1.990000E+2   -1.990000E+2   -2.388845E-4   -1.196864E-3   -7.685539E-5   3.489282E-6   -3.490490E-6   -7.685534E-5   7.693456E-5   1.774005E+2   2.673996E+2   
1.092326E+4   2.043841E+1   2.043841E+1   -1.490000E+2   -1.490000E+2   8.999910E+1   -1.490000E+2   -1.490000E+2   7.386554E-3   -7.020602E-3   -6.511358E-5   2.535989E-6   -2.537012E-6   -6.511354E-5   6.516294E-5   1.777696E+2   2.677687E+2   
1.095005E+4   2.042831E+1   2.042831E+1   -9.900000E+1   -9.900000E+1   8.999910E+1   -9.900000E+1   -9.900000E+1   1.485568E-2   -1.223678E-2   -5.385152E-5   1.263993E-6   -1.264838E-6   -5.385150E-5   5.386635E-5   1.786554E+2   2.686545E+2   
1.097679E+4   2.044619E+1   2.044619E+1   -4.900000E+1   -4.900000E+1   8.999910E+1   -4.800000E+1   -4.800000E+1   2.008220E-2   -1.963400E-2   -4.267751E-5   3.088666E-6   -3.089336E-6   -4.267746E-5   4.278913E-5   1.758606E+2   2.658597E+2   
1.100328E+4   2.044631E+1   2.044631E+1   0.000000E+0   0.000000E+0   8.999910E+1   0.000000E+0   0.000000E+0   2.696298E-2   -2.577980E-2   -3.135585E-5   2.869225E-6   -2.869717E-6   -3.135580E-5   3.148685E-5   1.747717E+2   2.647708E+2   
1.104161E+4   2.044540E+1   2.044540E+1   9.000000E+0   9.000000E+0   8.999910E+1   1.000000E+1   1.000000E+1   2.966443E-2   -2.652083E-2   -2.848414E-5   1.563417E-6   -1.563864E-6   -2.848411E-5   2.852701E-5   1.768583E+2   2.668574E+2   
1.106840E+4   2.042471E+1   2.042471E+1   1.900000E+1   1.900000E+1   8.999910E+1   2.000000E+1   2.000000E+1   3.071963E-2   -2.765005E-2   -2.647136E-5   1.674180E-6   -1.674595E-6   -2.647133E-5   2.652425E-5   1.763812E+2   2.663803E+2   
1.109525E+4   2.043099E+1   2.043099E+1   2.900000E+1   2.900000E+1   8.999910E+1   3.000000E+1   3.000000E+1   3.226476E-2   -2.936399E-2   -2.377027E-5   1.855832E-6   -1.856205E-6   -2.377024E-5   2.384260E-5   1.755358E+2   2.655349E+2   
1.112214E+4   2.042391E+1   2.042391E+1   3.900000E+1   3.900000E+1   8.999910E+1   4.000000E+1   4.000000E+1   3.224525E-2   -3.015012E-2   -2.268681E-5   2.471853E-6   -2.472209E-6   -2.268677E-5   2.282107E-5   1.737818E+2   2.637809E+2   
1.114895E+4   2.042159E+1   2.042159E+1   4.900000E+1   4.900000E+1   8.999910E+1   4.900000E+1   4.900000E+1   3.455853E-2   -3.107488E-2   -2.002172E-5   1.559938E-6   -1.560253E-6   -2.002170E-5   2.008240E-5   1.755450E+2   2.655441E+2   
1.117585E+4   2.040099E+1   2.040099E+1   5.900000E+1   5.900000E+1   8.999910E+1   6.000000E+1   6.000000E+1   3.624565E-2   -3.309260E-2   -1.697707E-5   1.861563E-6   -1.861830E-6   -1.697704E-5   1.707883E-5   1.737424E+2   2.637415E+2   
1.120273E+4   2.040649E+1   2.040649E+1   6.900000E+1   6.900000E+1   8.999910E+1   7.000000E+1   7.000000E+1   3.711098E-2   -3.318310E-2   -1.573286E-5   1.373710E-6   -1.373957E-6   -1.573284E-5   1.579272E-5   1.750099E+2   2.650090E+2   
1.122962E+4   2.041070E+1   2.041070E+1   7.900000E+1   7.900000E+1   8.999910E+1   7.900000E+1   7.900000E+1   3.790166E-2   -3.454787E-2   -1.381216E-5   1.828916E-6   -1.829133E-6   -1.381213E-5   1.393272E-5   1.724571E+2   2.624562E+2   
1.125642E+4   2.039300E+1   2.039300E+1   8.900000E+1   8.900000E+1   8.999910E+1   8.900000E+1   8.900000E+1   3.979875E-2   -3.697787E-2   -1.043368E-5   2.269675E-6   -2.269839E-6   -1.043364E-5   1.067769E-5   1.677274E+2   2.577265E+2   
1.128322E+4   2.039630E+1   2.039630E+1   9.900000E+1   9.900000E+1   8.999910E+1   9.900000E+1   9.900000E+1   4.130094E-2   -3.706378E-2   -8.767232E-6   1.336198E-6   -1.336336E-6   -8.767211E-6   8.868472E-6   1.713343E+2   2.613334E+2   
1.131018E+4   2.038439E+1   2.038439E+1   1.090000E+2   1.090000E+2   8.999910E+1   1.090000E+2   1.090000E+2   4.248651E-2   -3.812323E-2   -6.710545E-6   1.307331E-6   -1.307436E-6   -6.710524E-6   6.836704E-6   1.689759E+2   2.589750E+2   
1.133723E+4   2.037551E+1   2.037551E+1   1.190000E+2   1.190000E+2   8.999910E+1   1.190000E+2   1.190000E+2   4.324094E-2   -4.122083E-2   -3.682210E-6   3.011335E-6   -3.011393E-6   -3.682163E-6   4.756765E-6   1.407235E+2   2.307226E+2   
1.136422E+4   2.039001E+1   2.039001E+1   1.290000E+2   1.290000E+2   8.999910E+1   1.300000E+2   1.300000E+2   4.580748E-2   -4.158799E-2   -1.070497E-6   1.541274E-6   -1.541291E-6   -1.070472E-6   1.876563E-6   1.247820E+2   2.147811E+2   
1.139126E+4   2.037139E+1   2.037139E+1   1.390000E+2   1.390000E+2   8.999910E+1   1.400000E+2   1.400000E+2   4.631725E-2   -4.291099E-2   6.979752E-7   2.167200E-6   -2.167190E-6   6.980092E-7   2.276824E-6   7.214817E+1   1.621473E+2   
1.141829E+4   2.036459E+1   2.036459E+1   1.490000E+2   1.490000E+2   8.999910E+1   1.500000E+2   1.500000E+2   4.746293E-2   -4.365660E-2   2.534105E-6   1.945326E-6   -1.945286E-6   2.534135E-6   3.194680E-6   3.751194E+1   1.275110E+2   
1.144528E+4   2.036779E+1   2.036779E+1   1.590000E+2   1.590000E+2   8.999910E+1   1.600000E+2   1.600000E+2   4.944504E-2   -4.601925E-2   5.927720E-6   2.279651E-6   -2.279558E-6   5.927756E-6   6.350958E-6   2.103548E+1   1.110346E+2   
1.147234E+4   2.036431E+1   2.036431E+1   1.690000E+2   1.690000E+2   8.999910E+1   1.690000E+2   1.690000E+2   5.107094E-2   -4.640134E-2   7.798684E-6   1.463582E-6   -1.463459E-6   7.798707E-6   7.934831E-6   1.062908E+1   1.006282E+2   
1.149940E+4   2.035470E+1   2.035470E+1   1.790000E+2   1.790000E+2   8.999910E+1   1.800000E+2   1.800000E+2   5.167546E-2   -4.728802E-2   9.421856E-6   1.721796E-6   -1.721648E-6   9.421883E-6   9.577889E-6   1.035624E+1   1.003553E+2   
1.152638E+4   2.035500E+1   2.035500E+1   1.890000E+2   1.890000E+2   8.999910E+1   1.890000E+2   1.890000E+2   5.174795E-2   -4.758205E-2   1.020158E-5   1.922864E-6   -1.922704E-6   1.020161E-5   1.038122E-5   1.067427E+1   1.006734E+2   
1.155340E+4   2.035690E+1   2.035690E+1   1.990000E+2   1.990000E+2   8.999910E+1   1.990000E+2   1.990000E+2   5.432482E-2   -4.974968E-2   1.387165E-5   1.706896E-6   -1.706678E-6   1.387168E-5   1.397627E-5   7.014940E+0   9.701404E+1   
1.158045E+4   2.035821E+1   2.035821E+1   2.090000E+2   2.090000E+2   8.999910E+1   2.100000E+2   2.100000E+2   5.590438E-2   -4.905803E-2   1.517034E-5   1.777945E-7   -1.775562E-7   1.517035E-5   1.517138E-5   6.714684E-1   9.067057E+1   
1.160755E+4   2.035079E+1   2.035079E+1   2.190000E+2   2.190000E+2   8.999910E+1   2.190000E+2   2.190000E+2   5.797483E-2   -5.234786E-2   1.913477E-5   1.097860E-6   -1.097559E-6   1.913479E-5   1.916624E-5   3.283752E+0   9.328285E+1   
1.163462E+4   2.035070E+1   2.035070E+1   2.290000E+2   2.290000E+2   8.999910E+1   2.290000E+2   2.290000E+2   5.969301E-2   -5.518160E-2   2.264331E-5   1.946835E-6   -1.946479E-6   2.264334E-5   2.272685E-5   4.914112E+0   9.491321E+1   
1.166163E+4   2.035519E+1   2.035519E+1   2.390000E+2   2.390000E+2   8.999910E+1   2.400000E+2   2.400000E+2   5.958179E-2   -5.616730E-2   2.384996E-5   2.771875E-6   -2.771500E-6   2.385000E-5   2.401049E-5   6.629254E+0   9.662835E+1   
1.168863E+4   2.035800E+1   2.035800E+1   2.490000E+2   2.490000E+2   8.999910E+1   2.500000E+2   2.500000E+2   6.262146E-2   -5.589399E-2   2.632062E-5   5.177639E-7   -5.173504E-7   2.632063E-5   2.632572E-5   1.126944E+0   9.112604E+1   
1.171568E+4   2.036141E+1   2.036141E+1   2.590000E+2   2.590000E+2   8.999910E+1   2.600000E+2   2.600000E+2   6.364223E-2   -5.773682E-2   2.875137E-5   1.154306E-6   -1.153854E-6   2.875139E-5   2.877454E-5   2.299068E+0   9.229817E+1   
1.174273E+4   2.036160E+1   2.036160E+1   2.690000E+2   2.690000E+2   8.999910E+1   2.690000E+2   2.690000E+2   6.465959E-2   -5.719812E-2   2.964719E-5   1.133818E-7   -1.129161E-7   2.964719E-5   2.964741E-5   2.191192E-1   9.021822E+1   
1.176978E+4   2.037740E+1   2.037740E+1   2.790000E+2   2.790000E+2   8.999910E+1   2.790000E+2   2.790000E+2   6.572939E-2   -6.058488E-2   3.306470E-5   1.801680E-6   -1.801160E-6   3.306473E-5   3.311375E-5   3.118935E+0   9.311804E+1   
1.179689E+4   2.037411E+1   2.037411E+1   2.890000E+2   2.890000E+2   8.999910E+1   2.890000E+2   2.890000E+2   6.831172E-2   -5.899434E-2   3.441618E-5   -1.061124E-6   1.061665E-6   3.441616E-5   3.443253E-5   -1.765992E+0   8.823311E+1   
1.182394E+4   2.037869E+1   2.037869E+1   2.990000E+2   2.990000E+2   8.999910E+1   2.990000E+2   2.990000E+2   6.982394E-2   -6.178233E-2   3.775898E-5   -1.012496E-7   1.018427E-7   3.775898E-5   3.775912E-5   -1.536366E-1   8.984546E+1   
1.185098E+4   2.036590E+1   2.036590E+1   3.090000E+2   3.090000E+2   8.999910E+1   3.100000E+2   3.100000E+2   6.911126E-2   -6.154315E-2   3.780730E-5   2.801631E-7   -2.795693E-7   3.780730E-5   3.780834E-5   4.245707E-1   9.042367E+1   
1.187806E+4   2.036941E+1   2.036941E+1   3.190000E+2   3.190000E+2   8.999910E+1   3.190000E+2   3.190000E+2   7.198943E-2   -7.155708E-2   4.646579E-5   5.368062E-6   -5.367332E-6   4.646587E-5   4.677484E-5   6.590006E+0   9.658911E+1   
1.190515E+4   2.037731E+1   2.037731E+1   3.290000E+2   3.290000E+2   8.999910E+1   3.290000E+2   3.290000E+2   6.958688E-2   -6.110255E-2   3.901287E-5   -2.658526E-7   2.664655E-7   3.901287E-5   3.901378E-5   -3.904352E-1   8.960866E+1   
1.193223E+4   2.036370E+1   2.036370E+1   3.390000E+2   3.390000E+2   8.999910E+1   3.390000E+2   3.390000E+2   7.385084E-2   -7.409430E-2   5.049742E-5   5.958612E-6   -5.957819E-6   5.049752E-5   5.084776E-5   6.729688E+0   9.672879E+1   
1.195929E+4   2.035659E+1   2.035659E+1   3.490000E+2   3.490000E+2   8.999910E+1   3.490000E+2   3.490000E+2   7.578874E-2   -6.752713E-2   4.834362E-5   4.350552E-8   -4.274614E-8   4.834362E-5   4.834364E-5   5.156176E-2   9.005066E+1   
1.198629E+4   2.035021E+1   2.035021E+1   3.590000E+2   3.590000E+2   8.999910E+1   3.590000E+2   3.590000E+2   7.623176E-2   -6.364374E-2   4.685042E-5   -2.945745E-6   2.946481E-6   4.685038E-5   4.694294E-5   -3.597767E+0   8.640133E+1   
1.201329E+4   2.034670E+1   2.034670E+1   3.690000E+2   3.690000E+2   8.999910E+1   3.690000E+2   3.690000E+2   7.843200E-2   -7.076730E-2   5.333147E-5   5.853057E-7   -5.844680E-7   5.333148E-5   5.333469E-5   6.287882E-1   9.062789E+1   
1.204039E+4   2.033831E+1   2.033831E+1   3.790000E+2   3.790000E+2   8.999910E+1   3.790000E+2   3.790000E+2   7.898747E-2   -7.267138E-2   5.548952E-5   1.588148E-6   -1.587277E-6   5.548954E-5   5.551224E-5   1.639397E+0   9.163850E+1   
1.206739E+4   2.032360E+1   2.032360E+1   3.890000E+2   3.890000E+2   8.999910E+1   3.890000E+2   3.890000E+2   8.148204E-2   -8.719911E-2   6.674219E-5   1.012193E-5   -1.012088E-5   6.674235E-5   6.750536E-5   8.623603E+0   9.862270E+1   
1.209446E+4   2.033590E+1   2.033590E+1   3.990000E+2   3.990000E+2   8.999910E+1   4.000000E+2   4.000000E+2   8.194639E-2   -7.245501E-2   5.861327E-5   -5.152698E-7   5.161905E-7   5.861326E-5   5.861553E-5   -5.036748E-1   8.949543E+1   
1.212162E+4   2.033810E+1   2.033810E+1   4.090000E+2   4.090000E+2   8.999910E+1   4.090000E+2   4.090000E+2   8.344825E-2   -7.406204E-2   6.115835E-5   -3.837091E-7   3.846698E-7   6.115834E-5   6.115955E-5   -3.594705E-1   8.963963E+1   
1.214866E+4   2.033019E+1   2.033019E+1   4.190000E+2   4.190000E+2   8.999910E+1   4.190000E+2   4.190000E+2   8.454064E-2   -7.638721E-2   6.393495E-5   5.423017E-7   -5.412974E-7   6.393496E-5   6.393725E-5   4.859760E-1   9.048508E+1   
1.217571E+4   2.032049E+1   2.032049E+1   4.290000E+2   4.290000E+2   8.999910E+1   4.290000E+2   4.290000E+2   8.745024E-2   -8.061279E-2   6.909876E-5   1.542512E-6   -1.541427E-6   6.909878E-5   6.911597E-5   1.278818E+0   9.127792E+1   
1.220274E+4   2.031481E+1   2.031481E+1   4.390000E+2   4.390000E+2   8.999910E+1   4.390000E+2   4.390000E+2   8.825066E-2   -7.623942E-2   6.754133E-5   -2.039594E-6   2.040655E-6   6.754130E-5   6.757212E-5   -1.729676E+0   8.826942E+1   
1.222980E+4   2.031240E+1   2.031240E+1   4.490000E+2   4.490000E+2   8.999910E+1   4.490000E+2   4.490000E+2   8.892770E-2   -8.080477E-2   7.142496E-5   7.504091E-7   -7.492872E-7   7.142497E-5   7.142890E-5   6.019421E-1   9.060104E+1   
1.225690E+4   2.031350E+1   2.031350E+1   4.590000E+2   4.590000E+2   8.999910E+1   4.590000E+2   4.590000E+2   9.173802E-2   -8.283954E-2   7.516876E-5   2.788402E-7   -2.776595E-7   7.516876E-5   7.516928E-5   2.125390E-1   9.021164E+1   
1.228395E+4   2.031500E+1   2.031500E+1   4.680000E+2   4.680000E+2   8.999910E+1   4.690000E+2   4.690000E+2   9.266033E-2   -8.451572E-2   7.743082E-5   8.665726E-7   -8.653563E-7   7.743083E-5   7.743567E-5   6.412031E-1   9.064030E+1   
1.231100E+4   2.032110E+1   2.032110E+1   4.790000E+2   4.790000E+2   8.999910E+1   4.790000E+2   4.790000E+2   9.470950E-2   -8.302664E-2   7.848913E-5   -1.554506E-6   1.555739E-6   7.848911E-5   7.850452E-5   -1.134616E+0   8.886448E+1   
1.233805E+4   2.033611E+1   2.033611E+1   4.880000E+2   4.880000E+2   8.999910E+1   4.890000E+2   4.890000E+2   9.509530E-2   -8.553859E-2   8.090954E-5   -6.302656E-9   7.573580E-9   8.090954E-5   8.090954E-5   -4.463202E-3   8.999464E+1   
1.236503E+4   2.032549E+1   2.032549E+1   4.990000E+2   4.990000E+2   8.999910E+1   4.990000E+2   4.990000E+2   9.752958E-2   -8.838633E-2   8.490469E-5   3.550790E-7   -3.537454E-7   8.490470E-5   8.490543E-5   2.396147E-1   9.023871E+1   
1.239209E+4   2.033520E+1   2.033520E+1   5.090000E+2   5.090000E+2   8.999910E+1   5.090000E+2   5.090000E+2   9.821212E-2   -8.759865E-2   8.548426E-5   -6.234038E-7   6.247466E-7   8.548425E-5   8.548653E-5   -4.178287E-1   8.958127E+1   
1.241919E+4   2.034380E+1   2.034380E+1   5.190000E+2   5.190000E+2   8.999910E+1   5.190000E+2   5.190000E+2   9.976611E-2   -8.704472E-2   8.678991E-5   -2.042853E-6   2.044216E-6   8.678988E-5   8.681395E-5   -1.348374E+0   8.865073E+1   
1.244623E+4   2.033560E+1   2.033560E+1   5.280000E+2   5.280000E+2   8.999910E+1   5.290000E+2   5.290000E+2   1.012247E-1   -9.017856E-2   9.031066E-5   -8.025257E-7   8.039443E-7   9.031064E-5   9.031422E-5   -5.091329E-1   8.948997E+1   
1.247318E+4   2.034249E+1   2.034249E+1   5.380000E+2   5.380000E+2   8.999910E+1   5.390000E+2   5.390000E+2   1.040325E-1   -9.217129E-2   9.402679E-5   -1.301913E-6   1.303390E-6   9.402677E-5   9.403581E-5   -7.932779E-1   8.920582E+1   
1.250024E+4   2.033730E+1   2.033730E+1   5.480000E+2   5.480000E+2   8.999910E+1   5.490000E+2   5.490000E+2   1.032169E-1   -8.807851E-2   9.156409E-5   -3.564078E-6   3.565516E-6   9.156403E-5   9.163343E-5   -2.229079E+0   8.777002E+1   
1.252732E+4   2.033679E+1   2.033679E+1   5.580000E+2   5.580000E+2   8.999910E+1   5.590000E+2   5.590000E+2   1.066990E-1   -9.567660E-2   9.919395E-5   -5.897386E-7   5.912968E-7   9.919394E-5   9.919570E-5   -3.406371E-1   8.965846E+1   
1.255438E+4   2.036160E+1   2.036160E+1   5.680000E+2   5.680000E+2   8.999910E+1   5.690000E+2   5.690000E+2   1.084336E-1   -9.404855E-2   9.995647E-5   -2.890091E-6   2.891661E-6   9.995642E-5   9.999824E-5   -1.656160E+0   8.834294E+1   
1.258141E+4   2.033679E+1   2.033679E+1   5.780000E+2   5.780000E+2   8.999910E+1   5.790000E+2   5.790000E+2   1.085040E-1   -1.000875E-1   1.043458E-4   1.357703E-6   -1.356064E-6   1.043458E-4   1.043546E-4   7.454663E-1   9.074457E+1   
1.260874E+4   2.033792E+1   2.033792E+1   5.880000E+2   5.880000E+2   8.999910E+1   5.880000E+2   5.880000E+2   1.120784E-1   -9.914623E-2   1.066995E-4   -1.742608E-6   1.744284E-6   1.066995E-4   1.067137E-4   -9.356671E-1   8.906343E+1   
1.263604E+4   2.034969E+1   2.034969E+1   5.980000E+2   5.980000E+2   8.999910E+1   5.980000E+2   5.980000E+2   1.123664E-1   -9.922153E-2   1.075490E-4   -1.840076E-6   1.841765E-6   1.075489E-4   1.075647E-4   -9.801891E-1   8.901891E+1   
1.266330E+4   2.034850E+1   2.034850E+1   6.080000E+2   6.080000E+2   8.999910E+1   6.080000E+2   6.080000E+2   1.142530E-1   -1.046181E-1   1.127536E-4   6.942540E-7   -6.924829E-7   1.127536E-4   1.127557E-4   3.527809E-1   9.035188E+1   
1.269065E+4   2.035241E+1   2.035241E+1   6.180000E+2   6.180000E+2   8.999910E+1   6.180000E+2   6.180000E+2   1.166169E-1   -1.053537E-1   1.153966E-4   -3.809003E-7   3.827129E-7   1.153966E-4   1.153972E-4   -1.891208E-1   8.980998E+1   
1.271800E+4   2.035339E+1   2.035339E+1   6.280000E+2   6.280000E+2   8.999910E+1   6.280000E+2   6.280000E+2   1.164609E-1   -1.052848E-1   1.158606E-4   -2.713816E-7   2.732016E-7   1.158606E-4   1.158610E-4   -1.342043E-1   8.986490E+1   
1.274504E+4   2.033331E+1   2.033331E+1   6.380000E+2   6.380000E+2   8.999910E+1   6.390000E+2   6.390000E+2   1.183031E-1   -1.063092E-1   1.183950E-4   -7.760573E-7   7.779171E-7   1.183950E-4   1.183976E-4   -3.755578E-1   8.962354E+1   
1.277212E+4   2.032189E+1   2.032189E+1   6.480000E+2   6.480000E+2   8.999910E+1   6.480000E+2   6.480000E+2   1.204768E-1   -1.066752E-1   1.206217E-4   -1.984017E-6   1.985912E-6   1.206216E-4   1.206380E-4   -9.423311E-1   8.905677E+1   
1.279919E+4   2.033880E+1   2.033880E+1   6.580000E+2   6.580000E+2   8.999910E+1   6.580000E+2   6.580000E+2   1.224306E-1   -1.104035E-1   1.248402E-4   -6.695203E-7   6.714813E-7   1.248402E-4   1.248420E-4   -3.072754E-1   8.969182E+1   
1.282623E+4   2.034030E+1   2.034030E+1   6.680000E+2   6.680000E+2   8.999910E+1   6.680000E+2   6.680000E+2   1.246156E-1   -1.108270E-1   1.271710E-4   -1.839890E-6   1.841887E-6   1.271710E-4   1.271843E-4   -8.288883E-1   8.917021E+1   
1.285329E+4   2.031771E+1   2.031771E+1   6.780000E+2   6.780000E+2   8.999910E+1   6.780000E+2   6.780000E+2   1.253085E-1   -1.131367E-1   1.296714E-4   -6.472795E-7   6.493164E-7   1.296714E-4   1.296730E-4   -2.860005E-1   8.971310E+1   
1.288035E+4   2.033010E+1   2.033010E+1   6.880000E+2   6.880000E+2   8.999910E+1   6.880000E+2   6.880000E+2   1.287677E-1   -1.147333E-1   1.335775E-4   -1.877757E-6   1.879855E-6   1.335775E-4   1.335907E-4   -8.053783E-1   8.919372E+1   
1.290739E+4   2.036031E+1   2.036031E+1   6.980000E+2   6.980000E+2   8.999910E+1   6.980000E+2   6.980000E+2   1.319244E-1   -1.185140E-1   1.386314E-4   -1.362073E-6   1.364251E-6   1.386313E-4   1.386381E-4   -5.629211E-1   8.943618E+1   
1.293438E+4   2.033969E+1   2.033969E+1   7.080000E+2   7.080000E+2   8.999910E+1   7.080000E+2   7.080000E+2   1.323199E-1   -1.192949E-1   1.399886E-4   -1.037992E-6   1.040191E-6   1.399886E-4   1.399925E-4   -4.248307E-1   8.957427E+1   
1.296145E+4   2.034081E+1   2.034081E+1   7.180000E+2   7.180000E+2   8.999910E+1   7.180000E+2   7.180000E+2   1.333211E-1   -1.223044E-1   1.431273E-4   4.326267E-7   -4.303784E-7   1.431273E-4   1.431279E-4   1.731858E-1   9.017229E+1   
1.298878E+4   2.033300E+1   2.033300E+1   7.280000E+2   7.280000E+2   8.999910E+1   7.280000E+2   7.280000E+2   1.365863E-1   -1.222170E-1   1.458633E-4   -1.847402E-6   1.849694E-6   1.458632E-4   1.458750E-4   -7.256296E-1   8.927347E+1   
1.301633E+4   2.034399E+1   2.034399E+1   7.380000E+2   7.380000E+2   8.999910E+1   7.380000E+2   7.380000E+2   1.379724E-1   -1.249964E-1   1.491166E-4   -8.058989E-7   8.082412E-7   1.491166E-4   1.491188E-4   -3.096513E-1   8.968945E+1   
1.304357E+4   2.034710E+1   2.034710E+1   7.480000E+2   7.480000E+2   8.999910E+1   7.480000E+2   7.480000E+2   1.402320E-1   -1.255946E-1   1.516051E-4   -1.905327E-6   1.907709E-6   1.516051E-4   1.516171E-4   -7.200380E-1   8.927906E+1   
1.307111E+4   2.033679E+1   2.033679E+1   7.580000E+2   7.580000E+2   8.999910E+1   7.580000E+2   7.580000E+2   1.420142E-1   -1.301748E-1   1.562356E-4   1.274685E-7   -1.250144E-7   1.562356E-4   1.562356E-4   4.674611E-2   9.004585E+1   
1.309841E+4   2.034881E+1   2.034881E+1   7.680000E+2   7.680000E+2   8.999910E+1   7.680000E+2   7.680000E+2   1.442095E-1   -1.302915E-1   1.583837E-4   -1.265852E-6   1.268340E-6   1.583837E-4   1.583888E-4   -4.579160E-1   8.954118E+1   
1.312570E+4   2.035290E+1   2.035290E+1   7.780000E+2   7.780000E+2   8.999910E+1   7.780000E+2   7.780000E+2   1.458369E-1   -1.331996E-1   1.618776E-4   -3.015550E-7   3.040978E-7   1.618776E-4   1.618779E-4   -1.067338E-1   8.989237E+1   
1.315300E+4   2.035031E+1   2.035031E+1   7.880000E+2   7.880000E+2   8.999910E+1   7.880000E+2   7.880000E+2   1.467708E-1   -1.334403E-1   1.632604E-4   -7.314113E-7   7.339758E-7   1.632604E-4   1.632620E-4   -2.566851E-1   8.974241E+1   
1.318000E+4   2.035861E+1   2.035861E+1   7.980000E+2   7.980000E+2   8.999910E+1   7.980000E+2   7.980000E+2   1.495595E-1   -1.361390E-1   1.673999E-4   -7.209767E-7   7.236062E-7   1.673999E-4   1.674015E-4   -2.467663E-1   8.975233E+1   
1.320705E+4   2.035220E+1   2.035220E+1   8.080000E+2   8.080000E+2   8.999910E+1   8.080000E+2   8.080000E+2   1.513541E-1   -1.393587E-1   1.711981E-4   3.463535E-7   -3.436643E-7   1.711981E-4   1.711984E-4   1.159158E-1   9.011502E+1   
1.323408E+4   2.035531E+1   2.035531E+1   8.180000E+2   8.180000E+2   8.999910E+1   8.190000E+2   8.190000E+2   1.534267E-1   -1.393603E-1   1.732542E-4   -1.037715E-6   1.040437E-6   1.732541E-4   1.732573E-4   -3.431721E-1   8.965593E+1   
1.326105E+4   2.035150E+1   2.035150E+1   8.280000E+2   8.280000E+2   8.999910E+1   8.280000E+2   8.280000E+2   1.568853E-1   -1.418000E-1   1.776198E-4   -1.679804E-6   1.682594E-6   1.776198E-4   1.776278E-4   -5.418471E-1   8.945725E+1   
1.328832E+4   2.034350E+1   2.034350E+1   8.380000E+2   8.380000E+2   8.999910E+1   8.380000E+2   8.380000E+2   1.569710E-1   -1.430627E-1   1.790679E-4   -8.016819E-7   8.044947E-7   1.790679E-4   1.790697E-4   -2.565098E-1   8.974259E+1   
1.331534E+4   2.034850E+1   2.034850E+1   8.480000E+2   8.480000E+2   8.999910E+1   8.480000E+2   8.480000E+2   1.596544E-1   -1.459789E-1   1.832718E-4   -5.652031E-7   5.680819E-7   1.832718E-4   1.832726E-4   -1.766974E-1   8.982240E+1   
1.334263E+4   2.033651E+1   2.033651E+1   8.580000E+2   8.580000E+2   8.999910E+1   8.580000E+2   8.580000E+2   1.626179E-1   -1.483842E-1   1.873467E-4   -8.825942E-7   8.855371E-7   1.873467E-4   1.873488E-4   -2.699196E-1   8.972918E+1   
1.336968E+4   2.033361E+1   2.033361E+1   8.680000E+2   8.680000E+2   8.999910E+1   8.680000E+2   8.680000E+2   1.658124E-1   -1.519032E-1   1.922640E-4   -5.772157E-7   5.802358E-7   1.922640E-4   1.922649E-4   -1.720130E-1   8.982709E+1   
1.339691E+4   2.033370E+1   2.033370E+1   8.780000E+2   8.780000E+2   8.999910E+1   8.780000E+2   8.780000E+2   1.668612E-1   -1.554411E-1   1.957609E-4   1.231972E-6   -1.228897E-6   1.957609E-4   1.957648E-4   3.605718E-1   9.035967E+1   
1.342398E+4   2.032269E+1   2.032269E+1   8.880000E+2   8.880000E+2   8.999910E+1   8.880000E+2   8.880000E+2   1.710880E-1   -1.582760E-1   2.009446E-4   3.391610E-7   -3.360045E-7   2.009446E-4   2.009448E-4   9.670564E-2   9.009581E+1   
1.345128E+4   2.032519E+1   2.032519E+1   8.980000E+2   8.980000E+2   8.999910E+1   8.980000E+2   8.980000E+2   1.721108E-1   -1.600959E-1   2.033626E-4   9.581652E-7   -9.549708E-7   2.033626E-4   2.033648E-4   2.699534E-1   9.026905E+1   
1.347822E+4   2.031799E+1   2.031799E+1   9.080000E+2   9.080000E+2   8.999910E+1   9.080000E+2   9.080000E+2   1.771473E-1   -1.630655E-1   2.091699E-4   -4.023476E-7   4.056333E-7   2.091699E-4   2.091703E-4   -1.102109E-1   8.988889E+1   
1.350543E+4   2.031191E+1   2.031191E+1   9.180000E+2   9.180000E+2   8.999910E+1   9.180000E+2   9.180000E+2   1.789183E-1   -1.665117E-1   2.130921E-4   8.406751E-7   -8.373279E-7   2.130921E-4   2.130938E-4   2.260379E-1   9.022514E+1   
1.353249E+4   2.031411E+1   2.031411E+1   9.280000E+2   9.280000E+2   8.999910E+1   9.280000E+2   9.280000E+2   1.801782E-1   -1.737911E-1   2.190418E-4   5.134505E-6   -5.131064E-6   2.190419E-4   2.191020E-4   1.342810E+0   9.134191E+1   
1.355974E+4   2.032339E+1   2.032339E+1   9.380000E+2   9.380000E+2   8.999910E+1   9.380000E+2   9.380000E+2   1.817166E-1   -1.680547E-1   2.171347E-4   8.113327E-8   -7.772252E-8   2.171348E-4   2.171348E-4   2.140880E-2   9.002051E+1   
1.358680E+4   2.030001E+1   2.030001E+1   9.480000E+2   9.480000E+2   8.999910E+1   9.480000E+2   9.480000E+2   1.885363E-1   -1.779987E-1   2.284418E-4   2.386860E-6   -2.383271E-6   2.284419E-4   2.284543E-4   5.986294E-1   9.059773E+1   
1.361383E+4   2.029601E+1   2.029601E+1   9.580000E+2   9.580000E+2   8.999910E+1   9.590000E+2   9.590000E+2   1.978449E-1   -1.992546E-1   2.484611E-4   1.092410E-5   -1.092020E-5   2.484613E-4   2.487011E-4   2.517505E+0   9.251660E+1   
1.364115E+4   2.032339E+1   2.032339E+1   9.680000E+2   9.680000E+2   8.999910E+1   9.680000E+2   9.680000E+2   1.948255E-1   -1.850187E-1   2.381988E-4   3.054317E-6   -3.050576E-6   2.381988E-4   2.382184E-4   7.346381E-1   9.073374E+1   
1.366814E+4   2.031899E+1   2.031899E+1   9.780000E+2   9.780000E+2   8.999910E+1   9.780000E+2   9.780000E+2   2.008014E-1   -1.890326E-1   2.452784E-4   1.775663E-6   -1.771810E-6   2.452784E-4   2.452848E-4   4.147785E-1   9.041388E+1   
1.369546E+4   2.031240E+1   2.031240E+1   9.880000E+2   9.880000E+2   8.999910E+1   9.880000E+2   9.880000E+2   2.047524E-1   -1.953093E-1   2.524047E-4   3.494943E-6   -3.490978E-6   2.524048E-4   2.524289E-4   7.933000E-1   9.079240E+1   
1.372250E+4   2.030859E+1   2.030859E+1   9.980000E+2   9.980000E+2   8.999910E+1   9.990000E+2   9.990000E+2   2.075962E-1   -1.979280E-1   2.565927E-4   3.415733E-6   -3.411702E-6   2.565928E-4   2.566155E-4   7.626698E-1   9.076177E+1   
1.374996E+4   2.032479E+1   2.032479E+1   1.008000E+3   1.008000E+3   8.999910E+1   1.008000E+3   1.008000E+3   2.119071E-1   -2.031526E-1   2.632481E-4   4.140218E-6   -4.136083E-6   2.632482E-4   2.632807E-4   9.010415E-1   9.090014E+1   
1.377710E+4   2.033041E+1   2.033041E+1   1.018000E+3   1.018000E+3   8.999910E+1   1.019000E+3   1.019000E+3   2.149288E-1   -2.072266E-1   2.684541E-4   4.960869E-6   -4.956652E-6   2.684542E-4   2.684999E-4   1.058671E+0   9.105777E+1   
1.380459E+4   2.033080E+1   2.033080E+1   1.028000E+3   1.028000E+3   8.999910E+1   1.028000E+3   1.028000E+3   2.207348E-1   -2.108540E-1   2.751205E-4   3.523489E-6   -3.519168E-6   2.751205E-4   2.751430E-4   7.337515E-1   9.073285E+1   
1.383177E+4   2.034109E+1   2.034109E+1   1.038000E+3   1.038000E+3   8.999910E+1   1.039000E+3   1.039000E+3   2.260213E-1   -2.208256E-1   2.854824E-4   6.918534E-6   -6.914050E-6   2.854825E-4   2.855662E-4   1.388265E+0   9.138737E+1   
1.385926E+4   2.032821E+1   2.032821E+1   1.048000E+3   1.048000E+3   8.999910E+1   1.048000E+3   1.048000E+3   2.303669E-1   -2.233141E-1   2.904702E-4   5.694642E-6   -5.690079E-6   2.904703E-4   2.905260E-4   1.123135E+0   9.112223E+1   
1.388645E+4   2.031341E+1   2.031341E+1   1.058000E+3   1.058000E+3   8.999910E+1   1.058000E+3   1.058000E+3   2.342254E-1   -2.283279E-1   2.967543E-4   6.590051E-6   -6.585389E-6   2.967544E-4   2.968275E-4   1.272164E+0   9.127126E+1   
1.391408E+4   2.033209E+1   2.033209E+1   1.068000E+3   1.068000E+3   8.999910E+1   1.068000E+3   1.068000E+3   2.422182E-1   -2.385307E-1   3.090045E-4   8.262908E-6   -8.258055E-6   3.090046E-4   3.091149E-4   1.531748E+0   9.153085E+1   
1.394124E+4   2.032729E+1   2.032729E+1   1.078000E+3   1.078000E+3   8.999910E+1   1.078000E+3   1.078000E+3   2.466378E-1   -2.458429E-1   3.170834E-4   1.038493E-5   -1.037994E-5   3.170836E-4   3.172534E-4   1.875847E+0   9.187495E+1   
1.396872E+4   2.031280E+1   2.031280E+1   1.088000E+3   1.088000E+3   8.999910E+1   1.088000E+3   1.088000E+3   2.518080E-1   -2.585642E-1   3.290057E-4   1.578966E-5   -1.578449E-5   3.290059E-4   3.293844E-4   2.747633E+0   9.274673E+1   
1.399589E+4   2.030740E+1   2.030740E+1   1.098000E+3   1.098000E+3   8.999910E+1   1.098000E+3   1.098000E+3   2.565041E-1   -2.522083E-1   3.288234E-4   8.107145E-6   -8.101980E-6   3.288235E-4   3.289233E-4   1.412342E+0   9.141144E+1   
1.402334E+4   2.031149E+1   2.031149E+1   1.108000E+3   1.108000E+3   8.999910E+1   1.108000E+3   1.108000E+3   2.626698E-1   -2.618174E-1   3.394871E-4   1.063168E-5   -1.062635E-5   3.394872E-4   3.396535E-4   1.793739E+0   9.179284E+1   
1.405057E+4   2.030432E+1   2.030432E+1   1.118000E+3   1.118000E+3   8.999910E+1   1.119000E+3   1.119000E+3   2.670732E-1   -2.682909E-1   3.470980E-4   1.218005E-5   -1.217460E-5   3.470982E-4   3.473116E-4   2.009747E+0   9.200885E+1   
1.407783E+4   2.031161E+1   2.031161E+1   1.128000E+3   1.128000E+3   8.999910E+1   1.128000E+3   1.128000E+3   2.682202E-1   -2.749275E-1   3.525141E-4   1.609532E-5   -1.608978E-5   3.525144E-4   3.528814E-4   2.614232E+0   9.261333E+1   
1.410526E+4   2.030151E+1   2.030151E+1   1.138000E+3   1.138000E+3   8.999910E+1   1.139000E+3   1.139000E+3   2.724477E-1   -2.776354E-1   3.576808E-4   1.511764E-5   -1.511202E-5   3.576811E-4   3.580002E-4   2.420207E+0   9.241931E+1   
1.413244E+4   2.031750E+1   2.031750E+1   1.148000E+3   1.148000E+3   8.999910E+1   1.149000E+3   1.149000E+3   2.746545E-1   -2.786655E-1   3.604010E-4   1.435879E-5   -1.435312E-5   3.604012E-4   3.606869E-4   2.281523E+0   9.228062E+1   
1.415993E+4   2.031860E+1   2.031860E+1   1.158000E+3   1.158000E+3   8.999910E+1   1.159000E+3   1.159000E+3   2.760901E-1   -2.795369E-1   3.625084E-4   1.402396E-5   -1.401827E-5   3.625086E-4   3.627795E-4   2.215434E+0   9.221453E+1   
1.418712E+4   2.030880E+1   2.030880E+1   1.168000E+3   1.168000E+3   8.999910E+1   1.169000E+3   1.169000E+3   2.775736E-1   -2.825163E-1   3.659503E-4   1.513838E-5   -1.513263E-5   3.659505E-4   3.662633E-4   2.368822E+0   9.236792E+1   
1.421461E+4   2.031930E+1   2.031930E+1   1.178000E+3   1.178000E+3   8.999910E+1   1.179000E+3   1.179000E+3   2.759570E-1   -2.792086E-1   3.634381E-4   1.398474E-5   -1.397903E-5   3.634383E-4   3.637071E-4   2.203598E+0   9.220270E+1   
1.424180E+4   2.033550E+1   2.033550E+1   1.188000E+3   1.188000E+3   8.999910E+1   1.188000E+3   1.188000E+3   2.781140E-1   -2.814866E-1   3.668350E-4   1.413310E-5   -1.412734E-5   3.668353E-4   3.671072E-4   2.206351E+0   9.220545E+1   
1.426926E+4   2.032821E+1   2.032821E+1   1.198000E+3   1.198000E+3   8.999910E+1   1.199000E+3   1.199000E+3   2.767669E-1   -2.812919E-1   3.664874E-4   1.498646E-5   -1.498070E-5   3.664876E-4   3.667937E-4   2.341643E+0   9.234074E+1   
1.429647E+4   2.034591E+1   2.034591E+1   1.208000E+3   1.208000E+3   8.999910E+1   1.208000E+3   1.208000E+3   2.753565E-1   -2.812472E-1   3.660681E-4   1.597935E-5   -1.597359E-5   3.660683E-4   3.664166E-4   2.499448E+0   9.249855E+1   
1.432392E+4   2.033209E+1   2.033209E+1   1.218000E+3   1.218000E+3   8.999910E+1   1.218000E+3   1.218000E+3   2.760236E-1   -2.816981E-1   3.674026E-4   1.588273E-5   -1.587695E-5   3.674029E-4   3.677458E-4   2.475341E+0   9.247444E+1   
1.435116E+4   2.034271E+1   2.034271E+1   1.228000E+3   1.228000E+3   8.999910E+1   1.229000E+3   1.229000E+3   2.746256E-1   -2.785336E-1   3.651859E-4   1.468282E-5   -1.467709E-5   3.651862E-4   3.654810E-4   2.302419E+0   9.230152E+1   
1.437860E+4   2.034149E+1   2.034149E+1   1.238000E+3   1.238000E+3   8.999910E+1   1.239000E+3   1.239000E+3   2.741248E-1   -2.814080E-1   3.672385E-4   1.710183E-5   -1.709606E-5   3.672388E-4   3.676365E-4   2.666265E+0   9.266536E+1   
1.440580E+4   2.034551E+1   2.034551E+1   1.248000E+3   1.248000E+3   8.999910E+1   1.249000E+3   1.249000E+3   2.750845E-1   -2.774728E-1   3.660582E-4   1.371728E-5   -1.371153E-5   3.660584E-4   3.663151E-4   2.146038E+0   9.214514E+1   
1.443323E+4   2.033941E+1   2.033941E+1   1.258000E+3   1.258000E+3   8.999910E+1   1.258000E+3   1.258000E+3   2.729514E-1   -2.783290E-1   3.657131E-4   1.584582E-5   -1.584008E-5   3.657134E-4   3.660563E-4   2.480992E+0   9.248009E+1   
1.446048E+4   2.032849E+1   2.032849E+1   1.268000E+3   1.268000E+3   8.999910E+1   1.269000E+3   1.269000E+3   2.738844E-1   -2.776456E-1   3.665854E-4   1.477158E-5   -1.476582E-5   3.665856E-4   3.668829E-4   2.307489E+0   9.230659E+1   
1.448768E+4   2.032531E+1   2.032531E+1   1.278000E+3   1.278000E+3   8.999910E+1   1.279000E+3   1.279000E+3   2.722504E-1   -2.768991E-1   3.656443E-4   1.543129E-5   -1.542555E-5   3.656445E-4   3.659697E-4   2.416621E+0   9.241572E+1   
1.451511E+4   2.032900E+1   2.032900E+1   1.288000E+3   1.288000E+3   8.999910E+1   1.289000E+3   1.289000E+3   2.736671E-1   -2.763621E-1   3.668687E-4   1.411911E-5   -1.411335E-5   3.668689E-4   3.671403E-4   2.203967E+0   9.220307E+1   
1.454234E+4   2.032830E+1   2.032830E+1   1.298000E+3   1.298000E+3   8.999910E+1   1.299000E+3   1.299000E+3   2.740958E-1   -2.756787E-1   3.673433E-4   1.339024E-5   -1.338447E-5   3.673435E-4   3.675872E-4   2.087597E+0   9.208670E+1   
1.456979E+4   2.032281E+1   2.032281E+1   1.308000E+3   1.308000E+3   8.999910E+1   1.309000E+3   1.309000E+3   2.721569E-1   -2.770912E-1   3.675327E-4   1.578010E-5   -1.577433E-5   3.675330E-4   3.678713E-4   2.458498E+0   9.245760E+1   
1.459700E+4   2.033419E+1   2.033419E+1   1.318000E+3   1.318000E+3   8.999910E+1   1.319000E+3   1.319000E+3   2.721064E-1   -2.767272E-1   3.678848E-4   1.560884E-5   -1.560306E-5   3.678850E-4   3.682158E-4   2.429523E+0   9.242862E+1   
1.462442E+4   2.033041E+1   2.033041E+1   1.328000E+3   1.328000E+3   8.999910E+1   1.329000E+3   1.329000E+3   2.720116E-1   -2.761361E-1   3.680670E-4   1.530853E-5   -1.530275E-5   3.680673E-4   3.683852E-4   2.381655E+0   9.238076E+1   
1.465167E+4   2.031970E+1   2.031970E+1   1.338000E+3   1.338000E+3   8.999910E+1   1.339000E+3   1.339000E+3   2.710359E-1   -2.740520E-1   3.667387E-4   1.457016E-5   -1.456440E-5   3.667389E-4   3.670280E-4   2.275107E+0   9.227421E+1   
1.467912E+4   2.031729E+1   2.031729E+1   1.348000E+3   1.348000E+3   8.999910E+1   1.349000E+3   1.349000E+3   2.712395E-1   -2.744321E-1   3.677202E-4   1.474572E-5   -1.473994E-5   3.677204E-4   3.680157E-4   2.296352E+0   9.229545E+1   
1.470635E+4   2.030520E+1   2.030520E+1   1.358000E+3   1.358000E+3   8.999910E+1   1.359000E+3   1.359000E+3   2.705412E-1   -2.738292E-1   3.674923E-4   1.485638E-5   -1.485061E-5   3.674925E-4   3.677925E-4   2.315001E+0   9.231410E+1   
1.473379E+4   2.031100E+1   2.031100E+1   1.368000E+3   1.368000E+3   8.999910E+1   1.369000E+3   1.369000E+3   2.704893E-1   -2.756842E-1   3.692145E-4   1.624661E-5   -1.624082E-5   3.692148E-4   3.695718E-4   2.519571E+0   9.251867E+1   
1.476101E+4   2.030911E+1   2.030911E+1   1.378000E+3   1.378000E+3   8.999910E+1   1.379000E+3   1.379000E+3   2.697637E-1   -2.725413E-1   3.673989E-4   1.458993E-5   -1.458416E-5   3.673991E-4   3.676885E-4   2.274101E+0   9.227320E+1   
1.478847E+4   2.030740E+1   2.030740E+1   1.388000E+3   1.388000E+3   8.999910E+1   1.389000E+3   1.389000E+3   2.699504E-1   -2.746016E-1   3.694073E-4   1.595875E-5   -1.595295E-5   3.694076E-4   3.697519E-4   2.473695E+0   9.247279E+1   
1.481593E+4   2.031750E+1   2.031750E+1   1.399000E+3   1.399000E+3   8.999910E+1   1.399000E+3   1.399000E+3   2.686063E-1   -2.748665E-1   3.692846E-4   1.712833E-5   -1.712253E-5   3.692849E-4   3.696816E-4   2.655617E+0   9.265472E+1   
1.484362E+4   2.031710E+1   2.031710E+1   1.408000E+3   1.408000E+3   8.999910E+1   1.409000E+3   1.409000E+3   2.694384E-1   -2.725477E-1   3.690179E-4   1.496916E-5   -1.496337E-5   3.690182E-4   3.693214E-4   2.322922E+0   9.232202E+1   
1.487079E+4   2.032559E+1   2.032559E+1   1.418000E+3   1.418000E+3   8.999910E+1   1.419000E+3   1.419000E+3   2.675021E-1   -2.721111E-1   3.680665E-4   1.605671E-5   -1.605093E-5   3.680668E-4   3.684166E-4   2.497915E+0   9.249702E+1   
1.489845E+4   2.032400E+1   2.032400E+1   1.428000E+3   1.428000E+3   8.999910E+1   1.429000E+3   1.429000E+3   2.687223E-1   -2.722365E-1   3.695692E-4   1.534692E-5   -1.534111E-5   3.695694E-4   3.698877E-4   2.377927E+0   9.237703E+1   
1.492590E+4   2.034261E+1   2.034261E+1   1.439000E+3   1.439000E+3   8.999910E+1   1.439000E+3   1.439000E+3   2.687908E-1   -2.726505E-1   3.704814E-4   1.564010E-5   -1.563428E-5   3.704817E-4   3.708114E-4   2.417342E+0   9.241644E+1   
1.495303E+4   2.033099E+1   2.033099E+1   1.448000E+3   1.448000E+3   8.999910E+1   1.449000E+3   1.449000E+3   2.694260E-1   -2.727648E-1   3.715867E-4   1.532890E-5   -1.532307E-5   3.715869E-4   3.719027E-4   2.362258E+0   9.236136E+1   
1.498072E+4   2.032339E+1   2.032339E+1   1.459000E+3   1.459000E+3   8.999910E+1   1.459000E+3   1.459000E+3   2.699619E-1   -2.717721E-1   3.719417E-4   1.430808E-5   -1.430224E-5   3.719419E-4   3.722168E-4   2.203002E+0   9.220210E+1   
1.500820E+4   2.033669E+1   2.033669E+1   1.469000E+3   1.469000E+3   8.999910E+1   1.469000E+3   1.469000E+3   2.694598E-1   -2.735237E-1   3.732996E-4   1.593827E-5   -1.593241E-5   3.732999E-4   3.736397E-4   2.444796E+0   9.244390E+1   
1.503543E+4   2.032061E+1   2.032061E+1   1.479000E+3   1.479000E+3   8.999910E+1   1.479000E+3   1.479000E+3   2.695052E-1   -2.739042E-1   3.741757E-4   1.622395E-5   -1.621807E-5   3.741760E-4   3.745273E-4   2.482742E+0   9.248184E+1   
1.506263E+4   2.032220E+1   2.032220E+1   1.488000E+3   1.488000E+3   8.999910E+1   1.489000E+3   1.489000E+3   2.676560E-1   -2.716967E-1   3.721882E-4   1.600557E-5   -1.599972E-5   3.721885E-4   3.725322E-4   2.462428E+0   9.246153E+1   
1.509031E+4   2.032629E+1   2.032629E+1   1.499000E+3   1.499000E+3   8.999910E+1   1.499000E+3   1.499000E+3   2.682281E-1   -2.727984E-1   3.738616E-4   1.643260E-5   -1.642672E-5   3.738618E-4   3.742225E-4   2.516741E+0   9.251584E+1   
1.511779E+4   2.032989E+1   2.032989E+1   1.509000E+3   1.509000E+3   8.999910E+1   1.509000E+3   1.509000E+3   2.700484E-1   -2.722239E-1   3.753322E-4   1.481367E-5   -1.480777E-5   3.753325E-4   3.756244E-4   2.260185E+0   9.225929E+1   
1.514503E+4   2.032360E+1   2.032360E+1   1.519000E+3   1.519000E+3   8.999910E+1   1.519000E+3   1.519000E+3   2.667267E-1   -2.707869E-1   3.728379E-4   1.616013E-5   -1.615427E-5   3.728381E-4   3.731879E-4   2.481850E+0   9.248095E+1   
1.517247E+4   2.030709E+1   2.030709E+1   1.529000E+3   1.529000E+3   8.999910E+1   1.529000E+3   1.529000E+3   2.656718E-1   -2.695934E-1   3.720071E-4   1.610309E-5   -1.609724E-5   3.720073E-4   3.723554E-4   2.478617E+0   9.247772E+1   
1.520013E+4   2.032601E+1   2.032601E+1   1.539000E+3   1.539000E+3   8.999910E+1   1.539000E+3   1.539000E+3   2.667970E-1   -2.712167E-1   3.743718E-4   1.651275E-5   -1.650687E-5   3.743721E-4   3.747358E-4   2.525559E+0   9.252466E+1   
1.522753E+4   2.031301E+1   2.031301E+1   1.549000E+3   1.549000E+3   8.999910E+1   1.549000E+3   1.549000E+3   2.667273E-1   -2.706654E-1   3.745954E-4   1.622301E-5   -1.621713E-5   3.745956E-4   3.749465E-4   2.479821E+0   9.247892E+1   
1.525523E+4   2.031469E+1   2.031469E+1   1.559000E+3   1.559000E+3   8.999910E+1   1.559000E+3   1.559000E+3   2.676451E-1   -2.712556E-1   3.761834E-4   1.605019E-5   -1.604428E-5   3.761837E-4   3.765257E-4   2.443092E+0   9.244219E+1   
1.528272E+4   2.030941E+1   2.030941E+1   1.569000E+3   1.569000E+3   8.999910E+1   1.569000E+3   1.569000E+3   2.645243E-1   -2.687440E-1   3.731592E-4   1.650130E-5   -1.649544E-5   3.731594E-4   3.735238E-4   2.532001E+0   9.253110E+1   
1.531047E+4   2.030950E+1   2.030950E+1   1.579000E+3   1.579000E+3   8.999910E+1   1.579000E+3   1.579000E+3   2.671690E-1   -2.708428E-1   3.768320E-4   1.618979E-5   -1.618387E-5   3.768323E-4   3.771796E-4   2.460079E+0   9.245918E+1   
1.533793E+4   2.030251E+1   2.030251E+1   1.588000E+3   1.588000E+3   8.999910E+1   1.589000E+3   1.589000E+3   2.603920E-1   -2.575113E-1   3.646816E-4   1.157123E-5   -1.156550E-5   3.646818E-4   3.648652E-4   1.817367E+0   9.181647E+1   
1.536541E+4   2.030609E+1   2.030609E+1   1.599000E+3   1.599000E+3   8.999910E+1   1.599000E+3   1.599000E+3   2.752598E-1   -2.902343E-1   3.954360E-4   2.430634E-5   -2.430013E-5   3.954364E-4   3.961824E-4   3.517385E+0   9.351649E+1   
1.539306E+4   2.030779E+1   2.030779E+1   1.608000E+3   1.608000E+3   8.999910E+1   1.609000E+3   1.609000E+3   2.637074E-1   -2.670271E-1   3.739959E-4   1.605962E-5   -1.605375E-5   3.739961E-4   3.743405E-4   2.458807E+0   9.245791E+1   
1.542050E+4   2.031561E+1   2.031561E+1   1.619000E+3   1.619000E+3   8.999910E+1   1.619000E+3   1.619000E+3   2.615665E-1   -2.673674E-1   3.733880E-4   1.783577E-5   -1.782990E-5   3.733883E-4   3.738137E-4   2.734791E+0   9.273389E+1   
1.544820E+4   2.032360E+1   2.032360E+1   1.629000E+3   1.629000E+3   8.999910E+1   1.629000E+3   1.629000E+3   2.619705E-1   -2.650566E-1   3.728404E-4   1.597957E-5   -1.597371E-5   3.728407E-4   3.731827E-4   2.454137E+0   9.245324E+1   
1.547566E+4   2.032360E+1   2.032360E+1   1.638000E+3   1.638000E+3   8.999910E+1   1.639000E+3   1.639000E+3   2.628880E-1   -2.667975E-1   3.751392E-4   1.661616E-5   -1.661026E-5   3.751395E-4   3.755071E-4   2.536162E+0   9.253526E+1   
1.550339E+4   2.032919E+1   2.032919E+1   1.649000E+3   1.649000E+3   8.999910E+1   1.649000E+3   1.649000E+3   2.615951E-1   -2.657117E-1   3.742161E-4   1.680030E-5   -1.679442E-5   3.742164E-4   3.745931E-4   2.570547E+0   9.256965E+1   
1.553084E+4   2.033450E+1   2.033450E+1   1.659000E+3   1.659000E+3   8.999910E+1   1.659000E+3   1.659000E+3   2.613654E-1   -2.635255E-1   3.733227E-4   1.547189E-5   -1.546603E-5   3.733229E-4   3.736431E-4   2.373194E+0   9.237229E+1   
1.555831E+4   2.034341E+1   2.034341E+1   1.669000E+3   1.669000E+3   8.999910E+1   1.669000E+3   1.669000E+3   2.602996E-1   -2.648273E-1   3.740264E-4   1.717736E-5   -1.717149E-5   3.740267E-4   3.744206E-4   2.629492E+0   9.262859E+1   
1.558601E+4   2.032931E+1   2.032931E+1   1.679000E+3   1.679000E+3   8.999910E+1   1.679000E+3   1.679000E+3   2.587089E-1   -2.609589E-1   3.711850E-4   1.561142E-5   -1.560558E-5   3.711853E-4   3.715132E-4   2.408344E+0   9.240744E+1   
1.561366E+4   2.032989E+1   2.032989E+1   1.689000E+3   1.689000E+3   8.999910E+1   1.689000E+3   1.689000E+3   2.596669E-1   -2.639073E-1   3.742571E-4   1.706909E-5   -1.706321E-5   3.742574E-4   3.746461E-4   2.611332E+0   9.261043E+1   
1.564095E+4   2.033199E+1   2.033199E+1   1.699000E+3   1.699000E+3   8.999910E+1   1.699000E+3   1.699000E+3   2.584856E-1   -2.611282E-1   3.723620E-4   1.598480E-5   -1.597895E-5   3.723623E-4   3.727050E-4   2.458091E+0   9.245719E+1   
1.566810E+4   2.030520E+1   2.030520E+1   1.709000E+3   1.709000E+3   8.999910E+1   1.709000E+3   1.709000E+3   2.583340E-1   -2.607281E-1   3.726244E-4   1.585830E-5   -1.585245E-5   3.726246E-4   3.729617E-4   2.436947E+0   9.243605E+1   
1.569580E+4   2.031509E+1   2.031509E+1   1.719000E+3   1.719000E+3   8.999910E+1   1.719000E+3   1.719000E+3   2.584885E-1   -2.613919E-1   3.737484E-4   1.626744E-5   -1.626157E-5   3.737487E-4   3.741023E-4   2.492233E+0   9.249133E+1   
1.572303E+4   2.032321E+1   2.032321E+1   1.729000E+3   1.729000E+3   8.999910E+1   1.729000E+3   1.729000E+3   2.563681E-1   -2.609137E-1   3.726483E-4   1.745361E-5   -1.744776E-5   3.726486E-4   3.730568E-4   2.681585E+0   9.268068E+1   
1.575048E+4   2.031490E+1   2.031490E+1   1.739000E+3   1.739000E+3   8.999910E+1   1.739000E+3   1.739000E+3   2.571622E-1   -2.611677E-1   3.739460E-4   1.713028E-5   -1.712440E-5   3.739463E-4   3.743382E-4   2.622857E+0   9.262196E+1   
1.577793E+4   2.032049E+1   2.032049E+1   1.749000E+3   1.749000E+3   8.999910E+1   1.749000E+3   1.749000E+3   2.566289E-1   -2.577400E-1   3.720828E-4   1.513965E-5   -1.513380E-5   3.720830E-4   3.723906E-4   2.330018E+0   9.232912E+1   
1.580517E+4   2.031039E+1   2.031039E+1   1.759000E+3   1.759000E+3   8.999910E+1   1.759000E+3   1.759000E+3   2.534611E-1   -2.541786E-1   3.683785E-4   1.488513E-5   -1.487934E-5   3.683787E-4   3.686791E-4   2.313901E+0   9.231300E+1   
1.583241E+4   2.029971E+1   2.029971E+1   1.769000E+3   1.769000E+3   8.999910E+1   1.769000E+3   1.769000E+3   2.565483E-1   -2.720244E-1   3.820770E-4   2.534079E-5   -2.533478E-5   3.820774E-4   3.829164E-4   3.794515E+0   9.379361E+1   
1.585959E+4   2.028439E+1   2.028439E+1   1.779000E+3   1.779000E+3   8.999910E+1   1.779000E+3   1.779000E+3   2.511897E-1   -2.498492E-1   3.654087E-4   1.351734E-5   -1.351160E-5   3.654089E-4   3.656586E-4   2.118541E+0   9.211764E+1   
1.588674E+4   2.030599E+1   2.030599E+1   1.789000E+3   1.789000E+3   8.999910E+1   1.789000E+3   1.789000E+3   2.496245E-1   -2.621472E-1   3.725739E-4   2.330314E-5   -2.329729E-5   3.725742E-4   3.733019E-4   3.578980E+0   9.357808E+1   
1.591398E+4   2.030239E+1   2.030239E+1   1.799000E+3   1.799000E+3   8.999910E+1   1.799000E+3   1.799000E+3   2.543292E-1   -2.553806E-1   3.721435E-4   1.532589E-5   -1.532004E-5   3.721438E-4   3.724590E-4   2.358264E+0   9.235736E+1   
1.594139E+4   2.030181E+1   2.030181E+1   1.809000E+3   1.809000E+3   8.999910E+1   1.809000E+3   1.809000E+3   2.548864E-1   -2.580408E-1   3.747700E-4   1.685929E-5   -1.685340E-5   3.747702E-4   3.751490E-4   2.575755E+0   9.257485E+1   
1.596888E+4   2.029101E+1   2.029101E+1   1.819000E+3   1.819000E+3   8.999910E+1   1.819000E+3   1.819000E+3   2.538788E-1   -2.548416E-1   3.727313E-4   1.535882E-5   -1.535297E-5   3.727315E-4   3.730476E-4   2.359604E+0   9.235870E+1   
1.599658E+4   2.029641E+1   2.029641E+1   1.828000E+3   1.828000E+3   8.999910E+1   1.829000E+3   1.829000E+3   2.521800E-1   -2.538665E-1   3.716056E-4   1.590278E-5   -1.589694E-5   3.716059E-4   3.719457E-4   2.450465E+0   9.244956E+1   
1.602429E+4   2.029070E+1   2.029070E+1   1.839000E+3   1.839000E+3   8.999910E+1   1.839000E+3   1.839000E+3   2.515420E-1   -2.546414E-1   3.722693E-4   1.694044E-5   -1.693460E-5   3.722696E-4   3.726546E-4   2.605497E+0   9.260460E+1   
1.605169E+4   2.030169E+1   2.030169E+1   1.849000E+3   1.849000E+3   8.999910E+1   1.849000E+3   1.849000E+3   2.527207E-1   -2.538768E-1   3.731943E-4   1.563361E-5   -1.562775E-5   3.731946E-4   3.735217E-4   2.398795E+0   9.239789E+1   
1.607894E+4   2.030432E+1   2.030432E+1   1.859000E+3   1.859000E+3   8.999910E+1   1.859000E+3   1.859000E+3   2.502592E-1   -2.539377E-1   3.721997E-4   1.743589E-5   -1.743004E-5   3.722000E-4   3.726079E-4   2.682089E+0   9.268119E+1   
1.610659E+4   2.030050E+1   2.030050E+1   1.868000E+3   1.868000E+3   8.999910E+1   1.869000E+3   1.869000E+3   2.508022E-1   -2.543674E-1   3.734384E-4   1.741046E-5   -1.740460E-5   3.734387E-4   3.738440E-4   2.669314E+0   9.266841E+1   
1.613423E+4   2.032311E+1   2.032311E+1   1.879000E+3   1.879000E+3   8.999910E+1   1.879000E+3   1.879000E+3   2.511423E-1   -2.527678E-1   3.732877E-4   1.609885E-5   -1.609298E-5   3.732879E-4   3.736347E-4   2.469475E+0   9.246858E+1   
1.616167E+4   2.030432E+1   2.030432E+1   1.889000E+3   1.889000E+3   8.999910E+1   1.889000E+3   1.889000E+3   2.501404E-1   -2.522876E-1   3.729330E-4   1.650667E-5   -1.650081E-5   3.729333E-4   3.732981E-4   2.534358E+0   9.253346E+1   
1.618893E+4   2.032610E+1   2.032610E+1   1.899000E+3   1.899000E+3   8.999910E+1   1.899000E+3   1.899000E+3   2.490955E-1   -2.529686E-1   3.732671E-4   1.776104E-5   -1.775517E-5   3.732674E-4   3.736894E-4   2.724230E+0   9.272333E+1   
1.621660E+4   2.033489E+1   2.033489E+1   1.909000E+3   1.909000E+3   8.999910E+1   1.909000E+3   1.909000E+3   2.473782E-1   -2.515926E-1   3.718814E-4   1.803588E-5   -1.803004E-5   3.718817E-4   3.723185E-4   2.776614E+0   9.277571E+1   
1.624380E+4   2.032421E+1   2.032421E+1   1.919000E+3   1.919000E+3   8.999910E+1   1.920000E+3   1.920000E+3   2.470556E-1   -2.497824E-1   3.712193E-4   1.704151E-5   -1.703568E-5   3.712195E-4   3.716102E-4   2.628424E+0   9.262752E+1   
1.627100E+4   2.032189E+1   2.032189E+1   1.929000E+3   1.929000E+3   8.999910E+1   1.929000E+3   1.929000E+3   2.466389E-1   -2.488149E-1   3.708930E-4   1.669515E-5   -1.668932E-5   3.708933E-4   3.712686E-4   2.577337E+0   9.257644E+1   
1.629873E+4   2.032989E+1   2.032989E+1   1.939000E+3   1.939000E+3   8.999910E+1   1.939000E+3   1.939000E+3   2.463975E-1   -2.493231E-1   3.716566E-4   1.726981E-5   -1.726397E-5   3.716569E-4   3.720576E-4   2.660455E+0   9.265956E+1   
1.632596E+4   2.032000E+1   2.032000E+1   1.949000E+3   1.949000E+3   8.999910E+1   1.949000E+3   1.949000E+3   2.468012E-1   -2.483150E-1   3.719138E-4   1.633003E-5   -1.632419E-5   3.719140E-4   3.722721E-4   2.514134E+0   9.251323E+1   
1.635343E+4   2.030950E+1   2.030950E+1   1.959000E+3   1.959000E+3   8.999910E+1   1.959000E+3   1.959000E+3   2.470147E-1   -2.484185E-1   3.727310E-4   1.630412E-5   -1.629827E-5   3.727312E-4   3.730874E-4   2.504654E+0   9.250375E+1   
1.638066E+4   2.030120E+1   2.030120E+1   1.969000E+3   1.969000E+3   8.999910E+1   1.969000E+3   1.969000E+3   2.466277E-1   -2.495066E-1   3.737558E-4   1.738776E-5   -1.738189E-5   3.737561E-4   3.741600E-4   2.663578E+0   9.266268E+1   
1.640835E+4   2.030331E+1   2.030331E+1   1.979000E+3   1.979000E+3   8.999910E+1   1.979000E+3   1.979000E+3   2.447816E-1   -2.477918E-1   3.720747E-4   1.751378E-5   -1.750793E-5   3.720750E-4   3.724867E-4   2.694957E+0   9.269406E+1   
1.643560E+4   2.031750E+1   2.031750E+1   1.989000E+3   1.989000E+3   8.999910E+1   1.989000E+3   1.989000E+3   2.446248E-1   -2.461257E-1   3.715512E-4   1.650058E-5   -1.649475E-5   3.715515E-4   3.719174E-4   2.542834E+0   9.254193E+1   
1.646279E+4   2.030700E+1   2.030700E+1   1.999000E+3   1.999000E+3   8.999910E+1   1.999000E+3   1.999000E+3   2.437682E-1   -2.457926E-1   3.713844E-4   1.691095E-5   -1.690512E-5   3.713846E-4   3.717692E-4   2.607157E+0   9.260626E+1   
1.650370E+4   2.030001E+1   2.030001E+1   2.099000E+3   2.099000E+3   8.999910E+1   2.099000E+3   2.099000E+3   2.378204E-1   -2.404808E-1   3.702395E-4   1.780289E-5   -1.779707E-5   3.702398E-4   3.706673E-4   2.752935E+0   9.275204E+1   
1.653214E+4   2.031979E+1   2.031979E+1   2.199000E+3   2.199000E+3   8.999910E+1   2.199000E+3   2.199000E+3   2.333609E-1   -2.367428E-1   3.710604E-4   1.876780E-5   -1.876197E-5   3.710607E-4   3.715347E-4   2.895486E+0   9.289459E+1   
1.656054E+4   2.031771E+1   2.031771E+1   2.298000E+3   2.298000E+3   8.999910E+1   2.299000E+3   2.299000E+3   2.279741E-1   -2.302095E-1   3.695352E-4   1.841094E-5   -1.840513E-5   3.695355E-4   3.699935E-4   2.852225E+0   9.285133E+1   
1.658974E+4   2.030889E+1   2.030889E+1   2.398000E+3   2.398000E+3   8.999910E+1   2.399000E+3   2.399000E+3   2.225928E-1   -2.235993E-1   3.679661E-4   1.799624E-5   -1.799046E-5   3.679663E-4   3.684059E-4   2.799952E+0   9.279905E+1   
1.661839E+4   2.031030E+1   2.031030E+1   2.498000E+3   2.498000E+3   8.999910E+1   2.499000E+3   2.499000E+3   2.188752E-1   -2.203628E-1   3.695920E-4   1.879849E-5   -1.879269E-5   3.695923E-4   3.700698E-4   2.911716E+0   9.291082E+1   
1.664706E+4   2.032479E+1   2.032479E+1   2.598000E+3   2.598000E+3   8.999910E+1   2.598000E+3   2.598000E+3   2.124473E-1   -2.145326E-1   3.677453E-4   1.965446E-5   -1.964869E-5   3.677456E-4   3.682702E-4   3.059311E+0   9.305841E+1   
1.667622E+4   2.032571E+1   2.032571E+1   2.698000E+3   2.698000E+3   8.999910E+1   2.699000E+3   2.699000E+3   2.108571E-1   -2.097635E-1   3.699053E-4   1.790603E-5   -1.790022E-5   3.699055E-4   3.703384E-4   2.771357E+0   9.277046E+1   
1.670467E+4   2.033251E+1   2.033251E+1   2.798000E+3   2.798000E+3   8.999910E+1   2.799000E+3   2.799000E+3   2.025683E-1   -2.031987E-1   3.664237E-4   1.954292E-5   -1.953717E-5   3.664240E-4   3.669444E-4   3.052933E+0   9.305203E+1   
1.673304E+4   2.032809E+1   2.032809E+1   2.898000E+3   2.898000E+3   8.999910E+1   2.898000E+3   2.898000E+3   2.001176E-1   -2.001883E-1   3.689739E-4   1.961914E-5   -1.961334E-5   3.689742E-4   3.694951E-4   3.043674E+0   9.304277E+1   
1.676220E+4   2.032650E+1   2.032650E+1   2.998000E+3   2.998000E+3   8.999910E+1   2.999000E+3   2.999000E+3   1.950839E-1   -1.947365E-1   3.684136E-4   1.978261E-5   -1.977682E-5   3.684139E-4   3.689444E-4   3.073644E+0   9.307274E+1   
1.679063E+4   2.032260E+1   2.032260E+1   3.098000E+3   3.098000E+3   8.999910E+1   3.099000E+3   3.099000E+3   1.895169E-1   -1.891332E-1   3.673427E-4   2.020506E-5   -2.019929E-5   3.673430E-4   3.678979E-4   3.148284E+0   9.314738E+1   
1.681908E+4   2.032379E+1   2.032379E+1   3.198000E+3   3.198000E+3   8.999910E+1   3.199000E+3   3.199000E+3   1.829361E-1   -1.847643E-1   3.663580E-4   2.219980E-5   -2.219405E-5   3.663583E-4   3.670300E-4   3.467651E+0   9.346675E+1   
1.684827E+4   2.032791E+1   2.032791E+1   3.298000E+3   3.298000E+3   8.999910E+1   3.299000E+3   3.299000E+3   1.778616E-1   -1.759417E-1   3.636265E-4   2.001602E-5   -2.001031E-5   3.636268E-4   3.641770E-4   3.150697E+0   9.314980E+1   
1.687667E+4   2.032180E+1   2.032180E+1   3.398000E+3   3.398000E+3   8.999910E+1   3.399000E+3   3.399000E+3   1.738316E-1   -1.767607E-1   3.675500E-4   2.388747E-5   -2.388170E-5   3.675504E-4   3.683254E-4   3.718485E+0   9.371758E+1   
1.690508E+4   2.032049E+1   2.032049E+1   3.498000E+3   3.498000E+3   8.999910E+1   3.499000E+3   3.499000E+3   1.694823E-1   -1.694488E-1   3.662361E-4   2.226238E-5   -2.225663E-5   3.662364E-4   3.669121E-4   3.478557E+0   9.347766E+1   
1.693420E+4   2.030819E+1   2.030819E+1   3.599000E+3   3.599000E+3   8.999910E+1   3.599000E+3   3.599000E+3   1.694262E-1   -1.551214E-1   3.634527E-4   1.272120E-5   -1.271549E-5   3.634529E-4   3.636753E-4   2.004590E+0   9.200369E+1   
1.696265E+4   2.030630E+1   2.030630E+1   3.698000E+3   3.698000E+3   8.999910E+1   3.699000E+3   3.699000E+3   1.592470E-1   -1.589439E-1   3.651278E-4   2.297639E-5   -2.297065E-5   3.651282E-4   3.658500E-4   3.600702E+0   9.359980E+1   
1.699131E+4   2.030770E+1   2.030770E+1   3.799000E+3   3.799000E+3   8.999910E+1   3.799000E+3   3.799000E+3   1.552713E-1   -1.510098E-1   3.636788E-4   2.065421E-5   -2.064850E-5   3.636791E-4   3.642649E-4   3.250476E+0   9.324958E+1   
1.702048E+4   2.029260E+1   2.029260E+1   3.898000E+3   3.898000E+3   8.999910E+1   3.899000E+3   3.899000E+3   1.499102E-1   -1.467833E-1   3.635961E-4   2.190194E-5   -2.189622E-5   3.635965E-4   3.642552E-4   3.447160E+0   9.344626E+1   
1.704913E+4   2.030389E+1   2.030389E+1   3.999000E+3   3.999000E+3   8.999910E+1   3.999000E+3   3.999000E+3   1.436090E-1   -1.419962E-1   3.625395E-4   2.340835E-5   -2.340266E-5   3.625399E-4   3.632945E-4   3.694330E+0   9.369343E+1   
1.707748E+4   2.030901E+1   2.030901E+1   4.099000E+3   4.099000E+3   8.999910E+1   4.099000E+3   4.099000E+3   1.359824E-1   -1.358672E-1   3.597691E-4   2.489175E-5   -2.488610E-5   3.597695E-4   3.606292E-4   3.957879E+0   9.395698E+1   
1.710663E+4   2.029601E+1   2.029601E+1   4.198000E+3   4.198000E+3   8.999910E+1   4.199000E+3   4.199000E+3   1.330987E-1   -1.321553E-1   3.616580E-4   2.478039E-5   -2.477471E-5   3.616584E-4   3.625060E-4   3.919714E+0   9.391881E+1   
1.713504E+4   2.029510E+1   2.029510E+1   4.298000E+3   4.298000E+3   8.999910E+1   4.299000E+3   4.299000E+3   1.292790E-1   -1.253018E-1   3.609808E-4   2.310976E-5   -2.310409E-5   3.609812E-4   3.617198E-4   3.663040E+0   9.366214E+1   
1.716350E+4   2.028570E+1   2.028570E+1   4.398000E+3   4.398000E+3   8.999910E+1   4.399000E+3   4.399000E+3   1.236481E-1   -1.246546E-1   3.629298E-4   2.706206E-5   -2.705636E-5   3.629302E-4   3.639373E-4   4.264400E+0   9.426350E+1   
1.719311E+4   2.029620E+1   2.029620E+1   4.498000E+3   4.498000E+3   8.999910E+1   4.498000E+3   4.498000E+3   1.200762E-1   -1.144408E-1   3.602805E-4   2.285120E-5   -2.284554E-5   3.602809E-4   3.610044E-4   3.629188E+0   9.362829E+1   
1.722175E+4   2.030279E+1   2.030279E+1   4.598000E+3   4.598000E+3   8.999910E+1   4.598000E+3   4.598000E+3   1.113005E-1   -1.093361E-1   3.573761E-4   2.585319E-5   -2.584758E-5   3.573765E-4   3.583101E-4   4.137665E+0   9.413677E+1   
1.725065E+4   2.031371E+1   2.031371E+1   4.698000E+3   4.698000E+3   8.999910E+1   4.698000E+3   4.698000E+3   1.068342E-1   -1.059688E-1   3.584216E-4   2.708355E-5   -2.707792E-5   3.584220E-4   3.594434E-4   4.321252E+0   9.432035E+1   
1.728030E+4   2.030160E+1   2.030160E+1   4.798000E+3   4.798000E+3   8.999910E+1   4.798000E+3   4.798000E+3   1.025443E-1   -1.009626E-1   3.585720E-4   2.703873E-5   -2.703309E-5   3.585725E-4   3.595901E-4   4.312323E+0   9.431142E+1   
1.730920E+4   2.032330E+1   2.032330E+1   4.898000E+3   4.898000E+3   8.999910E+1   4.898000E+3   4.898000E+3   9.884519E-2   -9.694384E-2   3.597270E-4   2.727800E-5   -2.727235E-5   3.597275E-4   3.607598E-4   4.336424E+0   9.433552E+1   
1.733809E+4   2.032369E+1   2.032369E+1   4.997000E+3   4.997000E+3   8.999910E+1   4.998000E+3   4.998000E+3   9.223562E-2   -9.098209E-2   3.577388E-4   2.817254E-5   -2.816692E-5   3.577392E-4   3.588464E-4   4.502847E+0   9.450195E+1   
1.736780E+4   2.035760E+1   2.035760E+1   5.098000E+3   5.098000E+3   8.999910E+1   5.098000E+3   5.098000E+3   8.665686E-2   -8.622629E-2   3.571838E-4   2.919915E-5   -2.919354E-5   3.571842E-4   3.583753E-4   4.673439E+0   9.467254E+1   
1.739645E+4   2.034170E+1   2.034170E+1   5.198000E+3   5.198000E+3   8.999910E+1   5.198000E+3   5.198000E+3   7.980228E-2   -7.109179E-2   3.493640E-4   2.381290E-5   -2.380741E-5   3.493644E-4   3.501746E-4   3.899290E+0   9.389839E+1   
1.742530E+4   2.036041E+1   2.036041E+1   5.298000E+3   5.298000E+3   8.999910E+1   5.298000E+3   5.298000E+3   7.755508E-2   -8.100826E-2   3.600989E-4   3.284393E-5   -3.283828E-5   3.600994E-4   3.615936E-4   5.211420E+0   9.521052E+1   
1.745455E+4   2.035711E+1   2.035711E+1   5.398000E+3   5.398000E+3   8.999910E+1   5.398000E+3   5.398000E+3   8.200065E-2   -6.731476E-2   3.607118E-4   2.062147E-5   -2.061581E-5   3.607121E-4   3.613008E-4   3.271971E+0   9.327107E+1   
1.748321E+4   2.036309E+1   2.036309E+1   5.498000E+3   5.498000E+3   8.999910E+1   5.498000E+3   5.498000E+3   6.733820E-2   -6.446338E-2   3.552706E-4   2.929739E-5   -2.929181E-5   3.552711E-4   3.564766E-4   4.714228E+0   9.471333E+1   
1.751167E+4   2.036791E+1   2.036791E+1   5.598000E+3   5.598000E+3   8.999910E+1   5.598000E+3   5.598000E+3   6.062354E-2   -5.678981E-2   3.521545E-4   2.906105E-5   -2.905552E-5   3.521550E-4   3.533516E-4   4.717563E+0   9.471666E+1   
1.754085E+4   2.036611E+1   2.036611E+1   5.698000E+3   5.698000E+3   8.999910E+1   5.698000E+3   5.698000E+3   5.658593E-2   -5.441255E-2   3.540978E-4   3.068987E-5   -3.068431E-5   3.540983E-4   3.554253E-4   4.953481E+0   9.495258E+1   
1.756973E+4   2.036901E+1   2.036901E+1   5.798000E+3   5.798000E+3   8.999910E+1   5.798000E+3   5.798000E+3   5.137191E-2   -4.953336E-2   3.537100E-4   3.137634E-5   -3.137079E-5   3.537105E-4   3.550989E-4   5.069234E+0   9.506833E+1   
1.759863E+4   2.036819E+1   2.036819E+1   5.898000E+3   5.898000E+3   8.999910E+1   5.898000E+3   5.898000E+3   4.575264E-2   -4.333270E-2   3.522351E-4   3.141495E-5   -3.140942E-5   3.522356E-4   3.536333E-4   5.096579E+0   9.509568E+1   
1.762787E+4   2.037429E+1   2.037429E+1   5.998000E+3   5.998000E+3   8.999910E+1   5.998000E+3   5.998000E+3   4.262061E-2   -3.851142E-2   3.532727E-4   3.069589E-5   -3.069035E-5   3.532732E-4   3.546038E-4   4.965963E+0   9.496506E+1   
@@END Data.
@Time at end of measurement: 23:51:50
@Instrument  Changes:
@Emu Range: 20 uV
@END Instrument  Changes:
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   136.053        121.375        7.339          Coercive Field: Field at which M//H changes sign
Ms  emu                                 3.954E-4       -4.314E-4      4.134E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -3.136E-5      -3.212E-5      -3.837E-7      Remanent Magnetization: M at H=0        
S                                       0.079          0.074          0.077          Squareness: Mr/Ms                       
S*                                      0.330          0.122          0.226          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
