@Filename: c:\vsm-lv\Will\data\AJA1810b_Pt_CoFeB_Ir8\AJA1810b_Pt_CoFeB_Ir8_IP_fine.VHD
@Measurement Controlfilename: c:\vsm-lv\Will\Recipes\6_kOe inPlane loop (RT).VHC
@Signal Manipulation filename: C:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA1810b_Pt_CoFeB_Ir8
@Date: 18 November 2024    (2024-18-11)
@Time: 14:03:47
@Test ID: 
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 0.0009 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Applied Field to 5999.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Auto Range Signal to 9.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 4
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 10.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 6000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 100.0000 [Oe] Max Stepsize/Sweeprate = 100.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =   10.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To:  0.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =   10.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From:  0.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 10.0000 [Oe] Max Stepsize/Sweeprate = 10.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =   10.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -6000.0000 [Oe] Min Stepsize/Sweeprate = 100.0000 [Oe] Max Stepsize/Sweeprate = 100.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =   10.00 [sec] Up & Down = No
@Section 3 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 2 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.538
@Y Coils Correction Factor: 0.969
@Sample Shape Correction Factor: 0.928
@Coil Angle Alpha: 46.000
@Coil Angle Beta: -43.440
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
14999.000000   1.000000
15248.000000   0.999857
15498.000000   0.999857
15748.000000   0.999857
15999.000000   0.999857
16248.000000   0.999857
16498.000000   0.999857
16748.000000   0.999857
16998.000000   0.999710
17248.000000   0.999710
17498.000000   0.999857
17748.000000   0.999710
17998.000000   0.999857
18248.000000   0.999857
18498.000000   0.999857
18747.000000   0.999710
18997.000000   0.999857
19247.000000   0.999857
19498.000000   0.999857
19748.000000   0.999857
19998.000000   1.000000
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = Yes   Method = Angle Dependent Straight Line
Angular BG Signal array length = 25
Angle = 0.000000, Ofx = 5.511961E-6, Ofy = 7.255357E-5, Ofz = 0.000000E+0,Sx = -6.637759E-8, Sy = 3.436505E-9, Sz = 0.000000E+0
Angle = 15.000000, Ofx = 2.427508E-5, Ofy = 6.341217E-5, Ofz = 0.000000E+0,Sx = -6.122584E-8, Sy = 5.840215E-9, Sz = 0.000000E+0
Angle = 30.000000, Ofx = 3.849872E-5, Ofy = 5.614447E-5, Ofz = 0.000000E+0,Sx = -5.635123E-8, Sy = 5.018955E-9, Sz = 0.000000E+0
Angle = 45.000000, Ofx = 5.162249E-5, Ofy = 4.202634E-5, Ofz = 0.000000E+0,Sx = -5.340771E-8, Sy = 2.320584E-9, Sz = 0.000000E+0
Angle = 60.000000, Ofx = 5.888400E-5, Ofy = 2.821182E-5, Ofz = 0.000000E+0,Sx = -5.406333E-8, Sy = -1.140501E-9, Sz = 0.000000E+0
Angle = 75.000000, Ofx = 6.221306E-5, Ofy = 1.289058E-5, Ofz = 0.000000E+0,Sx = -5.702493E-8, Sy = -3.657483E-9, Sz = 0.000000E+0
Angle = 90.000000, Ofx = 6.528234E-5, Ofy = -3.469610E-6, Ofz = 0.000000E+0,Sx = -6.107239E-8, Sy = -4.959955E-9, Sz = 0.000000E+0
Angle = 105.000000, Ofx = 6.057411E-5, Ofy = -2.091353E-5, Ofz = 0.000000E+0,Sx = -6.580139E-8, Sy = -4.363769E-9, Sz = 0.000000E+0
Angle = 120.000000, Ofx = 5.108214E-5, Ofy = -3.497132E-5, Ofz = 0.000000E+0,Sx = -6.884862E-8, Sy = -3.031072E-9, Sz = 0.000000E+0
Angle = 135.000000, Ofx = 4.040625E-5, Ofy = -4.776267E-5, Ofz = 0.000000E+0,Sx = -7.079075E-8, Sy = -1.151461E-9, Sz = 0.000000E+0
Angle = 150.000000, Ofx = 2.815022E-5, Ofy = -5.275402E-5, Ofz = 0.000000E+0,Sx = -7.120194E-8, Sy = 2.952987E-10, Sz = 0.000000E+0
Angle = 165.000000, Ofx = 1.212763E-5, Ofy = -5.879891E-5, Ofz = 0.000000E+0,Sx = -6.933078E-8, Sy = 2.280793E-9, Sz = 0.000000E+0
Angle = 180.000000, Ofx = -1.503896E-6, Ofy = -5.933596E-5, Ofz = 0.000000E+0,Sx = -6.651357E-8, Sy = 4.300089E-9, Sz = 0.000000E+0
Angle = 195.000000, Ofx = -1.730048E-5, Ofy = -5.754707E-5, Ofz = 0.000000E+0,Sx = -6.233355E-8, Sy = 8.012817E-9, Sz = 0.000000E+0
Angle = 210.000000, Ofx = -3.045760E-5, Ofy = -5.052679E-5, Ofz = 0.000000E+0,Sx = -5.781798E-8, Sy = 6.626921E-9, Sz = 0.000000E+0
Angle = 225.000000, Ofx = -4.215979E-5, Ofy = -4.022672E-5, Ofz = 0.000000E+0,Sx = -5.424357E-8, Sy = 3.244164E-9, Sz = 0.000000E+0
Angle = 240.000000, Ofx = -4.971286E-5, Ofy = -2.831545E-5, Ofz = 0.000000E+0,Sx = -5.470668E-8, Sy = 5.438258E-11, Sz = 0.000000E+0
Angle = 255.000000, Ofx = -5.636146E-5, Ofy = -1.346311E-5, Ofz = 0.000000E+0,Sx = -5.652969E-8, Sy = -2.877288E-9, Sz = 0.000000E+0
Angle = 270.000000, Ofx = -5.608366E-5, Ofy = 3.241239E-6, Ofz = 0.000000E+0,Sx = -6.052403E-8, Sy = -4.749283E-9, Sz = 0.000000E+0
Angle = 285.000000, Ofx = -5.288340E-5, Ofy = 1.695085E-5, Ofz = 0.000000E+0,Sx = -6.466049E-8, Sy = -5.255801E-9, Sz = 0.000000E+0
Angle = 300.000000, Ofx = -4.592161E-5, Ofy = 3.148083E-5, Ofz = 0.000000E+0,Sx = -6.903811E-8, Sy = -4.123988E-9, Sz = 0.000000E+0
Angle = 315.000000, Ofx = -3.562648E-5, Ofy = 4.183753E-5, Ofz = 0.000000E+0,Sx = -7.195187E-8, Sy = -1.570295E-9, Sz = 0.000000E+0
Angle = 330.000000, Ofx = -2.158101E-5, Ofy = 4.883870E-5, Ofz = 0.000000E+0,Sx = -7.205703E-8, Sy = 1.349250E-9, Sz = 0.000000E+0
Angle = 345.000000, Ofx = -8.527411E-6, Ofy = 5.632367E-5, Ofz = 0.000000E+0,Sx = -7.020069E-8, Sy = 3.857333E-9, Sz = 0.000000E+0
Angle = 360.000000, Ofx = 4.810742E-6, Ofy = 5.580095E-5, Ofz = 0.000000E+0,Sx = -6.573828E-8, Sy = 6.096652E-9, Sz = 0.000000E+0
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 15 October 2024  12:22:06
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 4
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 14:03:47
@@Data
New Section: Section 0: 
3.724100E+1   1.982061E+1   1.982061E+1   5.998000E+3   5.998000E+3   9.000000E-4   5.999000E+3   5.999000E+3   -5.118286E-3   2.778158E-2   4.086663E-4   -1.137529E-4   4.086681E-4   -1.137465E-4   4.242027E-4   -1.555463E+1   -1.555373E+1   
6.562000E+1   1.982809E+1   1.982809E+1   5.898000E+3   5.898000E+3   9.000000E-4   5.899000E+3   5.899000E+3   1.564139E-3   3.332410E-2   4.105685E-4   -1.123742E-4   4.105703E-4   -1.123677E-4   4.256694E-4   -1.530719E+1   -1.530629E+1   
9.284700E+1   1.984600E+1   1.984600E+1   5.798000E+3   5.798000E+3   9.000000E-4   5.798000E+3   5.798000E+3   5.939152E-3   3.765691E-2   4.099507E-4   -1.117845E-4   4.099524E-4   -1.117780E-4   4.249180E-4   -1.525248E+1   -1.525158E+1   
1.209410E+2   1.985079E+1   1.985079E+1   5.697000E+3   5.697000E+3   9.000000E-4   5.698000E+3   5.698000E+3   1.055202E-2   4.279028E-2   4.101275E-4   -1.115342E-4   4.101292E-4   -1.115277E-4   4.250228E-4   -1.521366E+1   -1.521276E+1   
1.480510E+2   1.986169E+1   1.986169E+1   5.598000E+3   5.598000E+3   9.000000E-4   5.598000E+3   5.598000E+3   1.472245E-2   4.465761E-2   4.077000E-4   -1.095609E-4   4.077017E-4   -1.095545E-4   4.221645E-4   -1.504169E+1   -1.504079E+1   
1.752450E+2   1.985629E+1   1.985629E+1   5.498000E+3   5.498000E+3   9.000000E-4   5.498000E+3   5.498000E+3   1.977226E-2   4.975389E-2   4.081542E-4   -1.089961E-4   4.081559E-4   -1.089897E-4   4.224571E-4   -1.495172E+1   -1.495082E+1   
2.024450E+2   1.986071E+1   1.986071E+1   5.398000E+3   5.398000E+3   9.000000E-4   5.398000E+3   5.398000E+3   2.579336E-2   5.383450E-2   4.085689E-4   -1.071553E-4   4.085706E-4   -1.071489E-4   4.223871E-4   -1.469597E+1   -1.469507E+1   
2.303490E+2   1.986480E+1   1.986480E+1   5.298000E+3   5.298000E+3   9.000000E-4   5.298000E+3   5.298000E+3   3.048772E-2   5.832586E-2   4.083508E-4   -1.064539E-4   4.083525E-4   -1.064475E-4   4.219986E-4   -1.461136E+1   -1.461046E+1   
2.575530E+2   1.986010E+1   1.986010E+1   5.198000E+3   5.198000E+3   9.000000E-4   5.198000E+3   5.198000E+3   3.480390E-2   6.237663E-2   4.075601E-4   -1.057326E-4   4.075618E-4   -1.057262E-4   4.210518E-4   -1.454353E+1   -1.454263E+1   
2.847290E+2   1.985909E+1   1.985909E+1   5.098000E+3   5.098000E+3   9.000000E-4   5.098000E+3   5.098000E+3   4.137066E-2   6.423180E-2   4.067888E-4   -1.021525E-4   4.067904E-4   -1.021461E-4   4.194189E-4   -1.409658E+1   -1.409568E+1   
3.118760E+2   1.987240E+1   1.987240E+1   4.998000E+3   4.998000E+3   9.000000E-4   4.998000E+3   4.998000E+3   5.154667E-2   6.049178E-2   4.045898E-4   -9.270593E-5   4.045913E-4   -9.269958E-5   4.150751E-4   -1.290572E+1   -1.290482E+1   
3.390950E+2   1.985360E+1   1.985360E+1   4.898000E+3   4.898000E+3   9.000000E-4   4.898000E+3   4.898000E+3   4.426877E-2   7.380066E-2   4.022559E-4   -1.054439E-4   4.022576E-4   -1.054375E-4   4.158464E-4   -1.468854E+1   -1.468764E+1   
3.670160E+2   1.985119E+1   1.985119E+1   4.798000E+3   4.798000E+3   9.000000E-4   4.799000E+3   4.799000E+3   4.534980E-2   8.404409E-2   4.036393E-4   -1.107119E-4   4.036411E-4   -1.107056E-4   4.185473E-4   -1.533812E+1   -1.533722E+1   
3.941860E+2   1.986480E+1   1.986480E+1   4.698000E+3   4.698000E+3   9.000000E-4   4.699000E+3   4.699000E+3   5.948335E-2   7.716858E-2   4.019845E-4   -9.668647E-5   4.019860E-4   -9.668016E-5   4.134487E-4   -1.352406E+1   -1.352316E+1   
4.225260E+2   1.988671E+1   1.988671E+1   4.598000E+3   4.598000E+3   9.000000E-4   4.598000E+3   4.598000E+3   6.055833E-2   8.887743E-2   4.042615E-4   -1.028573E-4   4.042631E-4   -1.028509E-4   4.171414E-4   -1.427502E+1   -1.427412E+1   
4.496580E+2   1.988729E+1   1.988729E+1   4.498000E+3   4.498000E+3   9.000000E-4   4.498000E+3   4.498000E+3   6.588184E-2   9.040695E-2   4.023975E-4   -9.990569E-5   4.023990E-4   -9.989937E-5   4.146141E-4   -1.394325E+1   -1.394235E+1   
4.773380E+2   1.988079E+1   1.988079E+1   4.398000E+3   4.398000E+3   9.000000E-4   4.398000E+3   4.398000E+3   7.163594E-2   9.405544E-2   4.023228E-4   -9.797612E-5   4.023243E-4   -9.796980E-5   4.140808E-4   -1.368661E+1   -1.368571E+1   
5.054550E+2   1.990521E+1   1.990521E+1   4.298000E+3   4.298000E+3   9.000000E-4   4.299000E+3   4.299000E+3   7.621199E-2   9.864744E-2   4.021596E-4   -9.741928E-5   4.021612E-4   -9.741296E-5   4.137909E-4   -1.361704E+1   -1.361614E+1   
5.326180E+2   1.990099E+1   1.990099E+1   4.198000E+3   4.198000E+3   9.000000E-4   4.199000E+3   4.199000E+3   8.060734E-2   1.030798E-1   4.016923E-4   -9.688097E-5   4.016938E-4   -9.687466E-5   4.132102E-4   -1.355975E+1   -1.355885E+1   
5.598110E+2   1.988900E+1   1.988900E+1   4.098000E+3   4.098000E+3   9.000000E-4   4.099000E+3   4.099000E+3   8.510743E-2   1.055120E-1   3.998911E-4   -9.503675E-5   3.998926E-4   -9.503047E-5   4.110291E-4   -1.336871E+1   -1.336781E+1   
5.879290E+2   1.990429E+1   1.990429E+1   3.999000E+3   3.999000E+3   9.000000E-4   3.999000E+3   3.999000E+3   8.859032E-2   1.123246E-1   4.004639E-4   -9.657830E-5   4.004654E-4   -9.657201E-5   4.119450E-4   -1.355889E+1   -1.355799E+1   
6.158320E+2   1.991091E+1   1.991091E+1   3.898000E+3   3.898000E+3   9.000000E-4   3.899000E+3   3.899000E+3   9.157396E-2   1.135346E-1   3.967497E-4   -9.499095E-5   3.967512E-4   -9.498472E-5   4.079628E-4   -1.346446E+1   -1.346356E+1   
6.434700E+2   1.992480E+1   1.992480E+1   3.798000E+3   3.798000E+3   9.000000E-4   3.799000E+3   3.799000E+3   9.753954E-2   1.204484E-1   3.991183E-4   -9.493798E-5   3.991198E-4   -9.493171E-5   4.102543E-4   -1.338025E+1   -1.337935E+1   
6.716280E+2   1.990759E+1   1.990759E+1   3.698000E+3   3.698000E+3   9.000000E-4   3.699000E+3   3.699000E+3   1.010123E-1   1.232338E-1   3.968518E-4   -9.399773E-5   3.968533E-4   -9.399150E-5   4.078320E-4   -1.332542E+1   -1.332452E+1   
6.993130E+2   1.990859E+1   1.990859E+1   3.598000E+3   3.598000E+3   9.000000E-4   3.598000E+3   3.598000E+3   1.045794E-1   1.268152E-1   3.951443E-4   -9.348292E-5   3.951458E-4   -9.347672E-5   4.060518E-4   -1.331027E+1   -1.330937E+1   
7.271410E+2   1.991671E+1   1.991671E+1   3.498000E+3   3.498000E+3   9.000000E-4   3.498000E+3   3.498000E+3   1.105469E-1   1.330237E-1   3.970182E-4   -9.299292E-5   3.970197E-4   -9.298669E-5   4.077636E-4   -1.318265E+1   -1.318175E+1   
7.548290E+2   1.992730E+1   1.992730E+1   3.398000E+3   3.398000E+3   9.000000E-4   3.398000E+3   3.398000E+3   1.155959E-1   1.363995E-1   3.962619E-4   -9.136541E-5   3.962634E-4   -9.135919E-5   4.066585E-4   -1.298368E+1   -1.298278E+1   
7.829310E+2   1.992669E+1   1.992669E+1   3.298000E+3   3.298000E+3   9.000000E-4   3.298000E+3   3.298000E+3   1.202277E-1   1.378637E-1   3.938715E-4   -8.883510E-5   3.938729E-4   -8.882892E-5   4.037654E-4   -1.271001E+1   -1.270911E+1   
8.105360E+2   1.993020E+1   1.993020E+1   3.198000E+3   3.198000E+3   9.000000E-4   3.198000E+3   3.198000E+3   1.214057E-1   1.416984E-1   3.907489E-4   -9.007479E-5   3.907503E-4   -9.006865E-5   4.009964E-4   -1.298097E+1   -1.298007E+1   
8.381290E+2   1.996270E+1   1.996270E+1   3.098000E+3   3.098000E+3   9.000000E-4   3.098000E+3   3.098000E+3   1.262868E-1   1.494589E-1   3.929596E-4   -9.126887E-5   3.929610E-4   -9.126270E-5   4.034194E-4   -1.307570E+1   -1.307480E+1   
8.654220E+2   1.993621E+1   1.993621E+1   2.998000E+3   2.998000E+3   9.000000E-4   2.998000E+3   2.998000E+3   1.318883E-1   1.546970E-1   3.938967E-4   -9.042347E-5   3.938981E-4   -9.041728E-5   4.041423E-4   -1.292889E+1   -1.292799E+1   
8.932870E+2   1.996209E+1   1.996209E+1   2.897000E+3   2.897000E+3   9.000000E-4   2.898000E+3   2.898000E+3   1.336249E-1   1.571530E-1   3.901926E-4   -9.043841E-5   3.901940E-4   -9.043228E-5   4.005364E-4   -1.304953E+1   -1.304863E+1   
9.213960E+2   1.995889E+1   1.995889E+1   2.798000E+3   2.798000E+3   9.000000E-4   2.798000E+3   2.798000E+3   1.424140E-1   1.596676E-1   3.914287E-4   -8.578252E-5   3.914301E-4   -8.577637E-5   4.007182E-4   -1.236109E+1   -1.236019E+1   
9.488380E+2   1.997259E+1   1.997259E+1   2.697000E+3   2.697000E+3   9.000000E-4   2.698000E+3   2.698000E+3   1.448209E-1   1.629414E-1   3.887654E-4   -8.585542E-5   3.887668E-4   -8.584931E-5   3.981328E-4   -1.245338E+1   -1.245248E+1   
9.767320E+2   1.998708E+1   1.998708E+1   2.598000E+3   2.598000E+3   9.000000E-4   2.598000E+3   2.598000E+3   1.478074E-1   1.690313E-1   3.884851E-4   -8.728168E-5   3.884865E-4   -8.727557E-5   3.981693E-4   -1.266249E+1   -1.266159E+1   
1.004607E+3   1.999899E+1   1.999899E+1   2.498000E+3   2.498000E+3   9.000000E-4   2.498000E+3   2.498000E+3   1.513971E-1   1.677709E-1   3.834546E-4   -8.376328E-5   3.834559E-4   -8.375726E-5   3.924967E-4   -1.232234E+1   -1.232144E+1   
1.032022E+3   2.001449E+1   2.001449E+1   2.398000E+3   2.398000E+3   9.000000E-4   2.398000E+3   2.398000E+3   1.552357E-1   1.762933E-1   3.854768E-4   -8.612395E-5   3.854782E-4   -8.611789E-5   3.949807E-4   -1.259429E+1   -1.259339E+1   
1.059625E+3   2.002059E+1   2.002059E+1   2.298000E+3   2.298000E+3   9.000000E-4   2.298000E+3   2.298000E+3   1.597654E-1   1.730155E-1   3.796806E-4   -8.073154E-5   3.796819E-4   -8.072557E-5   3.881687E-4   -1.200403E+1   -1.200313E+1   
1.087227E+3   2.004351E+1   2.004351E+1   2.198000E+3   2.198000E+3   9.000000E-4   2.198000E+3   2.198000E+3   1.601840E-1   1.840471E-1   3.810918E-4   -8.692534E-5   3.810931E-4   -8.691936E-5   3.908797E-4   -1.284909E+1   -1.284819E+1   
1.114828E+3   2.005520E+1   2.005520E+1   2.098000E+3   2.098000E+3   9.000000E-4   2.098000E+3   2.098000E+3   1.603235E-1   1.780008E-1   3.702989E-4   -8.275234E-5   3.703002E-4   -8.274653E-5   3.794328E-4   -1.259716E+1   -1.259626E+1   
1.142823E+3   2.006350E+1   2.006350E+1   1.999000E+3   1.999000E+3   9.000000E-4   1.999000E+3   1.999000E+3   1.604741E-1   1.757253E-1   3.622318E-4   -8.090552E-5   3.622331E-4   -8.089983E-5   3.711571E-4   -1.259053E+1   -1.258963E+1   
1.181734E+3   2.008419E+1   2.008419E+1   1.948000E+3   1.948000E+3   9.000000E-4   1.948000E+3   1.948000E+3   1.601819E-1   1.745585E-1   3.578230E-4   -8.020423E-5   3.578243E-4   -8.019861E-5   3.667015E-4   -1.263375E+1   -1.263285E+1   
1.209138E+3   2.009280E+1   2.009280E+1   1.898000E+3   1.898000E+3   9.000000E-4   1.898000E+3   1.898000E+3   1.598753E-1   1.747760E-1   3.544442E-4   -8.037141E-5   3.544455E-4   -8.036584E-5   3.634422E-4   -1.277597E+1   -1.277507E+1   
1.236574E+3   2.009649E+1   2.009649E+1   1.848000E+3   1.848000E+3   9.000000E-4   1.848000E+3   1.848000E+3   1.593388E-1   1.707462E-1   3.479186E-4   -7.806749E-5   3.479198E-4   -7.806202E-5   3.565696E-4   -1.264681E+1   -1.264591E+1   
1.263988E+3   2.010620E+1   2.010620E+1   1.798000E+3   1.798000E+3   9.000000E-4   1.799000E+3   1.799000E+3   1.583718E-1   1.712767E-1   3.443674E-4   -7.887229E-5   3.443687E-4   -7.886688E-5   3.532843E-4   -1.290026E+1   -1.289936E+1   
1.291095E+3   2.010629E+1   2.010629E+1   1.748000E+3   1.748000E+3   9.000000E-4   1.748000E+3   1.748000E+3   1.572071E-1   1.681505E-1   3.379746E-4   -7.754258E-5   3.379758E-4   -7.753727E-5   3.467559E-4   -1.292192E+1   -1.292102E+1   
1.318200E+3   2.011611E+1   2.011611E+1   1.698000E+3   1.698000E+3   9.000000E-4   1.698000E+3   1.698000E+3   1.571213E-1   1.614658E-1   3.298951E-4   -7.329725E-5   3.298962E-4   -7.329206E-5   3.379397E-4   -1.252669E+1   -1.252579E+1   
1.345625E+3   2.011660E+1   2.011660E+1   1.648000E+3   1.648000E+3   9.000000E-4   1.648000E+3   1.648000E+3   1.559587E-1   1.626815E-1   3.266235E-4   -7.465260E-5   3.266247E-4   -7.464747E-5   3.350462E-4   -1.287430E+1   -1.287340E+1   
1.372736E+3   2.013250E+1   2.013250E+1   1.598000E+3   1.598000E+3   9.000000E-4   1.599000E+3   1.599000E+3   1.553838E-1   1.591823E-1   3.205108E-4   -7.270566E-5   3.205120E-4   -7.270063E-5   3.286538E-4   -1.278086E+1   -1.277996E+1   
1.400188E+3   2.012341E+1   2.012341E+1   1.548000E+3   1.548000E+3   9.000000E-4   1.548000E+3   1.548000E+3   1.555728E-1   1.607213E-1   3.183393E-4   -7.335525E-5   3.183404E-4   -7.335025E-5   3.266816E-4   -1.297622E+1   -1.297532E+1   
1.427589E+3   2.013009E+1   2.013009E+1   1.498000E+3   1.498000E+3   9.000000E-4   1.499000E+3   1.499000E+3   1.519879E-1   1.527291E-1   3.069758E-4   -7.064080E-5   3.069769E-4   -7.063598E-5   3.149988E-4   -1.295921E+1   -1.295831E+1   
1.455010E+3   2.013119E+1   2.013119E+1   1.448000E+3   1.448000E+3   9.000000E-4   1.448000E+3   1.448000E+3   1.480101E-1   1.379081E-1   2.904043E-4   -6.396195E-5   2.904053E-4   -6.395738E-5   2.973647E-4   -1.242116E+1   -1.242026E+1   
1.482416E+3   2.014031E+1   2.014031E+1   1.398000E+3   1.398000E+3   9.000000E-4   1.398000E+3   1.398000E+3   1.498462E-1   1.429645E-1   2.919169E-4   -6.568925E-5   2.919179E-4   -6.568466E-5   2.992166E-4   -1.268187E+1   -1.268097E+1   
1.509786E+3   2.013790E+1   2.013790E+1   1.348000E+3   1.348000E+3   9.000000E-4   1.348000E+3   1.348000E+3   1.476472E-1   1.486778E-1   2.910884E-4   -7.051555E-5   2.910895E-4   -7.051098E-5   2.995077E-4   -1.361745E+1   -1.361655E+1   
1.537224E+3   2.013409E+1   2.013409E+1   1.298000E+3   1.298000E+3   9.000000E-4   1.298000E+3   1.298000E+3   1.472686E-1   1.484051E-1   2.873147E-4   -7.042789E-5   2.873158E-4   -7.042338E-5   2.958206E-4   -1.377303E+1   -1.377213E+1   
1.564595E+3   2.012710E+1   2.012710E+1   1.248000E+3   1.248000E+3   9.000000E-4   1.248000E+3   1.248000E+3   1.429725E-1   1.492668E-1   2.816175E-4   -7.365587E-5   2.816186E-4   -7.365144E-5   2.910903E-4   -1.465715E+1   -1.465625E+1   
1.592019E+3   2.014190E+1   2.014190E+1   1.198000E+3   1.198000E+3   9.000000E-4   1.198000E+3   1.198000E+3   1.444047E-1   1.380708E-1   2.714198E-4   -6.560967E-5   2.714209E-4   -6.560540E-5   2.792371E-4   -1.358929E+1   -1.358839E+1   
1.619419E+3   2.014431E+1   2.014431E+1   1.148000E+3   1.148000E+3   9.000000E-4   1.148000E+3   1.148000E+3   1.448989E-1   1.494939E-1   2.764777E-4   -7.216680E-5   2.764789E-4   -7.216245E-5   2.857411E-4   -1.462906E+1   -1.462816E+1   
1.646839E+3   2.014810E+1   2.014810E+1   1.098000E+3   1.098000E+3   9.000000E-4   1.098000E+3   1.098000E+3   1.407920E-1   1.318252E-1   2.578802E-4   -6.381780E-5   2.578812E-4   -6.381375E-5   2.656594E-4   -1.389977E+1   -1.389887E+1   
1.674219E+3   2.016290E+1   2.016290E+1   1.048000E+3   1.048000E+3   9.000000E-4   1.048000E+3   1.048000E+3   1.396500E-1   1.330004E-1   2.545946E-4   -6.513438E-5   2.545956E-4   -6.513038E-5   2.627944E-4   -1.435050E+1   -1.434960E+1   
1.701497E+3   2.017639E+1   2.017639E+1   9.980000E+2   9.980000E+2   9.000000E-4   9.980000E+2   9.980000E+2   1.360147E-1   1.267792E-1   2.443752E-4   -6.354460E-5   2.443762E-4   -6.354076E-5   2.525018E-4   -1.457576E+1   -1.457486E+1   
1.728436E+3   2.018029E+1   2.018029E+1   9.470000E+2   9.470000E+2   9.000000E-4   9.480000E+2   9.480000E+2   1.317619E-1   1.246697E-1   2.366185E-4   -6.490761E-5   2.366195E-4   -6.490390E-5   2.453595E-4   -1.533967E+1   -1.533877E+1   
1.755368E+3   2.018499E+1   2.018499E+1   8.970000E+2   8.970000E+2   9.000000E-4   8.980000E+2   8.980000E+2   1.322105E-1   1.235741E-1   2.328408E-4   -6.375937E-5   2.328418E-4   -6.375571E-5   2.414127E-4   -1.531404E+1   -1.531314E+1   
1.782319E+3   2.019790E+1   2.019790E+1   8.470000E+2   8.470000E+2   9.000000E-4   8.480000E+2   8.480000E+2   1.281604E-1   1.212854E-1   2.250989E-4   -6.487633E-5   2.250999E-4   -6.487280E-5   2.342615E-4   -1.607765E+1   -1.607675E+1   
1.809353E+3   2.019061E+1   2.019061E+1   7.980000E+2   7.980000E+2   9.000000E-4   7.980000E+2   7.980000E+2   1.257547E-1   1.127993E-1   2.141410E-4   -6.106632E-5   2.141419E-4   -6.106296E-5   2.226779E-4   -1.591649E+1   -1.591559E+1   
1.836308E+3   2.019799E+1   2.019799E+1   7.470000E+2   7.470000E+2   9.000000E-4   7.480000E+2   7.480000E+2   1.228121E-1   1.077456E-1   2.052239E-4   -5.973559E-5   2.052248E-4   -5.973236E-5   2.137409E-4   -1.622897E+1   -1.622807E+1   
1.863272E+3   2.020281E+1   2.020281E+1   6.970000E+2   6.970000E+2   9.000000E-4   6.980000E+2   6.980000E+2   1.193517E-1   1.063531E-1   1.985219E-4   -6.101277E-5   1.985229E-4   -6.100965E-5   2.076861E-4   -1.708403E+1   -1.708313E+1   
1.890297E+3   2.020150E+1   2.020150E+1   6.480000E+2   6.480000E+2   9.000000E-4   6.480000E+2   6.480000E+2   1.117157E-1   1.022841E-1   1.870370E-4   -6.342306E-5   1.870380E-4   -6.342012E-5   1.974976E-4   -1.873147E+1   -1.873057E+1   
1.917236E+3   2.021441E+1   2.021441E+1   5.980000E+2   5.980000E+2   9.000000E-4   5.980000E+2   5.980000E+2   1.120131E-1   9.357642E-2   1.778010E-4   -5.767194E-5   1.778019E-4   -5.766914E-5   1.869204E-4   -1.797111E+1   -1.797021E+1   
1.944177E+3   2.020580E+1   2.020580E+1   5.480000E+2   5.480000E+2   9.000000E-4   5.480000E+2   5.480000E+2   1.025016E-1   9.670746E-2   1.700767E-4   -6.578315E-5   1.700777E-4   -6.578047E-5   1.823554E-4   -2.114573E+1   -2.114483E+1   
1.971076E+3   2.019711E+1   2.019711E+1   4.980000E+2   4.980000E+2   9.000000E-4   4.980000E+2   4.980000E+2   1.066837E-1   8.615666E-2   1.622431E-4   -5.630026E-5   1.622440E-4   -5.629771E-5   1.717339E-4   -1.913737E+1   -1.913647E+1   
1.998025E+3   2.020480E+1   2.020480E+1   4.480000E+2   4.480000E+2   9.000000E-4   4.480000E+2   4.480000E+2   9.928650E-2   7.609782E-2   1.467116E-4   -5.484980E-5   1.467125E-4   -5.484750E-5   1.566295E-4   -2.049882E+1   -2.049792E+1   
2.024981E+3   2.021389E+1   2.021389E+1   3.980000E+2   3.980000E+2   9.000000E-4   3.990000E+2   3.990000E+2   9.523161E-2   7.645547E-2   1.408939E-4   -5.760876E-5   1.408948E-4   -5.760655E-5   1.522165E-4   -2.223870E+1   -2.223780E+1   
2.051880E+3   2.021011E+1   2.021011E+1   3.480000E+2   3.480000E+2   9.000000E-4   3.480000E+2   3.480000E+2   8.751910E-2   6.918104E-2   1.270352E-4   -5.808589E-5   1.270361E-4   -5.808389E-5   1.396850E-4   -2.457189E+1   -2.457099E+1   
2.078848E+3   2.020059E+1   2.020059E+1   2.980000E+2   2.980000E+2   9.000000E-4   2.980000E+2   2.980000E+2   8.202000E-2   6.428864E-2   1.164556E-4   -5.856110E-5   1.164566E-4   -5.855927E-5   1.303508E-4   -2.669608E+1   -2.669518E+1   
2.105765E+3   2.021011E+1   2.021011E+1   2.480000E+2   2.480000E+2   9.000000E-4   2.490000E+2   2.490000E+2   7.354387E-2   6.127622E-2   1.051965E-4   -6.218844E-5   1.051975E-4   -6.218679E-5   1.222036E-4   -3.059006E+1   -3.058916E+1   
2.132685E+3   2.019991E+1   2.019991E+1   1.980000E+2   1.980000E+2   9.000000E-4   1.990000E+2   1.990000E+2   6.666239E-2   5.015067E-2   8.927319E-5   -5.973458E-5   8.927412E-5   -5.973318E-5   1.074147E-4   -3.378732E+1   -3.378642E+1   
2.159648E+3   2.019921E+1   2.019921E+1   1.480000E+2   1.480000E+2   9.000000E-4   1.490000E+2   1.490000E+2   5.892776E-2   3.642179E-2   7.092636E-5   -5.624144E-5   7.092724E-5   -5.624032E-5   9.051877E-5   -3.841285E+1   -3.841195E+1   
2.186553E+3   2.020641E+1   2.020641E+1   9.800000E+1   9.800000E+1   9.000000E-4   9.900000E+1   9.900000E+1   4.632489E-2   2.309830E-2   4.948280E-5   -5.624801E-5   4.948369E-5   -5.624723E-5   7.491586E-5   -4.866109E+1   -4.866019E+1   
2.213374E+3   2.021041E+1   2.021041E+1   4.900000E+1   4.900000E+1   9.000000E-4   4.900000E+1   4.900000E+1   3.185295E-2   9.653980E-3   2.665590E-5   -5.742739E-5   2.665680E-5   -5.742698E-5   6.331226E-5   -6.510083E+1   -6.509993E+1   
2.239846E+3   2.020089E+1   2.020089E+1   0.000000E+0   0.000000E+0   9.000000E-4   0.000000E+0   0.000000E+0   1.249182E-2   -9.983211E-3   -3.856192E-6   -5.804658E-5   -3.855281E-6   -5.804664E-5   5.817452E-5   -9.380073E+1   -9.379983E+1   
2.278124E+3   2.021261E+1   2.021261E+1   -9.000000E+0   -9.000000E+0   9.000000E-4   -9.000000E+0   -9.000000E+0   6.239357E-3   -1.067503E-2   -9.283506E-6   -6.176122E-5   -9.282536E-6   -6.176137E-5   6.245504E-5   -9.854830E+1   -9.854740E+1   
2.304771E+3   2.022421E+1   2.022421E+1   -1.900000E+1   -1.900000E+1   9.000000E-4   -1.900000E+1   -1.900000E+1   3.205604E-3   -1.695658E-2   -1.647229E-5   -5.987005E-5   -1.647135E-5   -5.987030E-5   6.209476E-5   -1.053834E+2   -1.053825E+2   
2.331501E+3   2.022610E+1   2.022610E+1   -2.900000E+1   -2.900000E+1   9.000000E-4   -2.900000E+1   -2.900000E+1   4.006816E-4   -2.206581E-2   -2.267766E-5   -5.855057E-5   -2.267674E-5   -5.855093E-5   6.278890E-5   -1.111723E+2   -1.111714E+2   
2.358175E+3   2.022021E+1   2.022021E+1   -3.900000E+1   -3.900000E+1   9.000000E-4   -3.900000E+1   -3.900000E+1   -3.540165E-3   -2.341822E-2   -2.703011E-5   -6.031073E-5   -2.702917E-5   -6.031116E-5   6.609093E-5   -1.141410E+2   -1.141401E+2   
2.384836E+3   2.022170E+1   2.022170E+1   -4.900000E+1   -4.900000E+1   9.000000E-4   -4.900000E+1   -4.900000E+1   -8.726017E-3   -2.686011E-2   -3.371688E-5   -6.161067E-5   -3.371591E-5   -6.161120E-5   7.023320E-5   -1.186900E+2   -1.186891E+2   
2.411484E+3   2.021761E+1   2.021761E+1   -6.000000E+1   -6.000000E+1   9.000000E-4   -5.900000E+1   -5.900000E+1   -1.109202E-2   -3.104656E-2   -3.896839E-5   -6.056847E-5   -3.896744E-5   -6.056909E-5   7.202136E-5   -1.227563E+2   -1.227554E+2   
2.438156E+3   2.023391E+1   2.023391E+1   -7.000000E+1   -7.000000E+1   9.000000E-4   -6.900000E+1   -6.900000E+1   -1.318623E-2   -3.615119E-2   -4.467683E-5   -5.877748E-5   -4.467590E-5   -5.877819E-5   7.382961E-5   -1.272385E+2   -1.272376E+2   
2.464832E+3   2.022390E+1   2.022390E+1   -7.900000E+1   -7.900000E+1   9.000000E-4   -7.900000E+1   -7.900000E+1   -1.732908E-2   -3.495938E-2   -4.738035E-5   -6.224465E-5   -4.737938E-5   -6.224540E-5   7.822592E-5   -1.272782E+2   -1.272773E+2   
2.491501E+3   2.023239E+1   2.023239E+1   -9.000000E+1   -9.000000E+1   9.000000E-4   -8.900000E+1   -8.900000E+1   -2.035461E-2   -3.908015E-2   -5.304384E-5   -6.168322E-5   -5.304287E-5   -6.168406E-5   8.135398E-5   -1.306935E+2   -1.306926E+2   
2.518174E+3   2.022851E+1   2.022851E+1   -9.900000E+1   -9.900000E+1   9.000000E-4   -9.900000E+1   -9.900000E+1   -2.344307E-2   -3.502288E-2   -5.299975E-5   -6.621734E-5   -5.299871E-5   -6.621817E-5   8.481574E-5   -1.286735E+2   -1.286726E+2   
2.544925E+3   2.021719E+1   2.021719E+1   -1.100000E+2   -1.100000E+2   9.000000E-4   -1.090000E+2   -1.090000E+2   -2.261167E-2   -5.174746E-2   -6.484769E-5   -5.529327E-5   -6.484682E-5   -5.529429E-5   8.522071E-5   -1.395470E+2   -1.395461E+2   
2.571728E+3   2.023480E+1   2.023480E+1   -1.200000E+2   -1.200000E+2   9.000000E-4   -1.190000E+2   -1.190000E+2   -2.545211E-2   -5.090694E-2   -6.689353E-5   -5.767409E-5   -6.689262E-5   -5.767514E-5   8.832352E-5   -1.392328E+2   -1.392319E+2   
2.598577E+3   2.022451E+1   2.022451E+1   -1.300000E+2   -1.300000E+2   9.000000E-4   -1.290000E+2   -1.290000E+2   -2.777546E-2   -5.354031E-2   -7.102320E-5   -5.756313E-5   -7.102230E-5   -5.756424E-5   9.142105E-5   -1.409758E+2   -1.409749E+2   
2.625369E+3   2.022549E+1   2.022549E+1   -1.400000E+2   -1.400000E+2   9.000000E-4   -1.390000E+2   -1.390000E+2   -3.214240E-2   -4.350696E-2   -6.766451E-5   -6.664341E-5   -6.766347E-5   -6.664447E-5   9.497278E-5   -1.354356E+2   -1.354347E+2   
2.652193E+3   2.021551E+1   2.021551E+1   -1.500000E+2   -1.500000E+2   9.000000E-4   -1.490000E+2   -1.490000E+2   -3.274862E-2   -5.551171E-2   -7.719185E-5   -5.959542E-5   -7.719091E-5   -5.959663E-5   9.752023E-5   -1.423303E+2   -1.423294E+2   
2.678956E+3   2.021240E+1   2.021240E+1   -1.600000E+2   -1.600000E+2   9.000000E-4   -1.590000E+2   -1.590000E+2   -3.512114E-2   -5.481275E-2   -7.901219E-5   -6.157647E-5   -7.901122E-5   -6.157771E-5   1.001728E-4   -1.420697E+2   -1.420688E+2   
2.705789E+3   2.022729E+1   2.022729E+1   -1.700000E+2   -1.700000E+2   9.000000E-4   -1.690000E+2   -1.690000E+2   -3.643593E-2   -5.810626E-2   -8.290550E-5   -6.038444E-5   -8.290455E-5   -6.038574E-5   1.025651E-4   -1.439322E+2   -1.439313E+2   
2.732570E+3   2.022689E+1   2.022689E+1   -1.800000E+2   -1.800000E+2   9.000000E-4   -1.790000E+2   -1.790000E+2   -3.752888E-2   -6.319980E-2   -8.791058E-5   -5.793203E-5   -8.790967E-5   -5.793341E-5   1.052824E-4   -1.466156E+2   -1.466147E+2   
2.759371E+3   2.021981E+1   2.021981E+1   -1.890000E+2   -1.890000E+2   9.000000E-4   -1.890000E+2   -1.890000E+2   -4.027713E-2   -5.608613E-2   -8.548073E-5   -6.412775E-5   -8.547972E-5   -6.412909E-5   1.068612E-4   -1.431227E+2   -1.431218E+2   
2.786164E+3   2.022650E+1   2.022650E+1   -1.990000E+2   -1.990000E+2   9.000000E-4   -1.990000E+2   -1.990000E+2   -4.151634E-2   -6.606975E-2   -9.402641E-5   -5.875119E-5   -9.402549E-5   -5.875267E-5   1.108723E-4   -1.480013E+2   -1.480004E+2   
2.812963E+3   2.023062E+1   2.023062E+1   -2.100000E+2   -2.100000E+2   9.000000E-4   -2.090000E+2   -2.090000E+2   -4.482814E-2   -5.463729E-2   -8.895081E-5   -6.799180E-5   -8.894974E-5   -6.799320E-5   1.119604E-4   -1.426066E+2   -1.426057E+2   
2.839772E+3   2.022799E+1   2.022799E+1   -2.200000E+2   -2.200000E+2   9.000000E-4   -2.190000E+2   -2.190000E+2   -4.677185E-2   -5.868430E-2   -9.381091E-5   -6.675391E-5   -9.380986E-5   -6.675538E-5   1.151372E-4   -1.445651E+2   -1.445642E+2   
2.866581E+3   2.024389E+1   2.024389E+1   -2.300000E+2   -2.300000E+2   9.000000E-4   -2.290000E+2   -2.290000E+2   -4.533168E-2   -7.119618E-2   -1.022733E-4   -5.802674E-5   -1.022724E-4   -5.802834E-5   1.175880E-4   -1.504308E+2   -1.504299E+2   
2.893371E+3   2.025021E+1   2.025021E+1   -2.390000E+2   -2.390000E+2   9.000000E-4   -2.390000E+2   -2.390000E+2   -4.705812E-2   -7.602263E-2   -1.075307E-4   -5.616219E-5   -1.075298E-4   -5.616388E-5   1.213138E-4   -1.524224E+2   -1.524215E+2   
2.920188E+3   2.025109E+1   2.025109E+1   -2.500000E+2   -2.500000E+2   9.000000E-4   -2.490000E+2   -2.490000E+2   -4.691690E-2   -7.270917E-2   -1.057661E-4   -5.808108E-5   -1.057652E-4   -5.808274E-5   1.206643E-4   -1.512268E+2   -1.512259E+2   
2.946981E+3   2.026000E+1   2.026000E+1   -2.590000E+2   -2.590000E+2   9.000000E-4   -2.590000E+2   -2.590000E+2   -5.225955E-2   -6.906220E-2   -1.075765E-4   -6.386617E-5   -1.075755E-4   -6.386786E-5   1.251063E-4   -1.493032E+2   -1.493023E+2   
2.973795E+3   2.025451E+1   2.025451E+1   -2.690000E+2   -2.690000E+2   9.000000E-4   -2.690000E+2   -2.690000E+2   -5.213525E-2   -7.642226E-2   -1.133299E-4   -5.920077E-5   -1.133290E-4   -5.920255E-5   1.278609E-4   -1.524185E+2   -1.524176E+2   
3.000601E+3   2.025640E+1   2.025640E+1   -2.800000E+2   -2.800000E+2   9.000000E-4   -2.800000E+2   -2.800000E+2   -5.123698E-2   -8.204749E-2   -1.173921E-4   -5.508737E-5   -1.173912E-4   -5.508921E-5   1.296747E-4   -1.548612E+2   -1.548603E+2   
3.027347E+3   2.025759E+1   2.025759E+1   -2.900000E+2   -2.900000E+2   9.000000E-4   -2.890000E+2   -2.890000E+2   -5.304905E-2   -8.000140E-2   -1.178093E-4   -5.753024E-5   -1.178084E-4   -5.753209E-5   1.311059E-4   -1.539722E+2   -1.539713E+2   
3.054189E+3   2.025939E+1   2.025939E+1   -3.000000E+2   -3.000000E+2   9.000000E-4   -2.990000E+2   -2.990000E+2   -5.454803E-2   -8.189086E-2   -1.208432E-4   -5.732876E-5   -1.208423E-4   -5.733066E-5   1.337522E-4   -1.546200E+2   -1.546191E+2   
3.080984E+3   2.026251E+1   2.026251E+1   -3.100000E+2   -3.100000E+2   9.000000E-4   -3.090000E+2   -3.090000E+2   -5.524519E-2   -8.238417E-2   -1.223382E-4   -5.745486E-5   -1.223373E-4   -5.745678E-5   1.351580E-4   -1.548434E+2   -1.548425E+2   
3.107791E+3   2.027560E+1   2.027560E+1   -3.190000E+2   -3.190000E+2   9.000000E-4   -3.190000E+2   -3.190000E+2   -5.539599E-2   -8.288770E-2   -1.234608E-4   -5.720999E-5   -1.234599E-4   -5.721193E-5   1.360719E-4   -1.551377E+2   -1.551368E+2   
3.134584E+3   2.028091E+1   2.028091E+1   -3.300000E+2   -3.300000E+2   9.000000E-4   -3.290000E+2   -3.290000E+2   -5.527885E-2   -7.944914E-2   -1.216250E-4   -5.922227E-5   -1.216241E-4   -5.922418E-5   1.352772E-4   -1.540374E+2   -1.540365E+2   
3.161390E+3   2.029479E+1   2.029479E+1   -3.400000E+2   -3.400000E+2   9.000000E-4   -3.390000E+2   -3.390000E+2   -5.707427E-2   -8.214287E-2   -1.254304E-4   -5.872165E-5   -1.254295E-4   -5.872362E-5   1.384956E-4   -1.549128E+2   -1.549119E+2   
3.188191E+3   2.029931E+1   2.029931E+1   -3.500000E+2   -3.500000E+2   9.000000E-4   -3.490000E+2   -3.490000E+2   -5.758633E-2   -8.478721E-2   -1.283096E-4   -5.739501E-5   -1.283086E-4   -5.739702E-5   1.405615E-4   -1.559002E+2   -1.558993E+2   
3.214984E+3   2.029659E+1   2.029659E+1   -3.590000E+2   -3.590000E+2   9.000000E-4   -3.590000E+2   -3.590000E+2   -5.831607E-2   -8.673470E-2   -1.308498E-4   -5.664426E-5   -1.308489E-4   -5.664631E-5   1.425842E-4   -1.565924E+2   -1.565915E+2   
3.241793E+3   2.029339E+1   2.029339E+1   -3.690000E+2   -3.690000E+2   9.000000E-4   -3.690000E+2   -3.690000E+2   -6.038819E-2   -8.626957E-2   -1.326259E-4   -5.828030E-5   -1.326250E-4   -5.828239E-5   1.448663E-4   -1.562777E+2   -1.562768E+2   
3.268608E+3   2.028121E+1   2.028121E+1   -3.790000E+2   -3.790000E+2   9.000000E-4   -3.790000E+2   -3.790000E+2   -6.175080E-2   -9.000369E-2   -1.368623E-4   -5.684792E-5   -1.368614E-4   -5.685007E-5   1.481991E-4   -1.574437E+2   -1.574428E+2   
3.295394E+3   2.028710E+1   2.028710E+1   -3.890000E+2   -3.890000E+2   9.000000E-4   -3.890000E+2   -3.890000E+2   -6.298422E-2   -8.972411E-2   -1.381863E-4   -5.780955E-5   -1.381854E-4   -5.781172E-5   1.497912E-4   -1.572982E+2   -1.572973E+2   
3.322201E+3   2.026541E+1   2.026541E+1   -3.990000E+2   -3.990000E+2   9.000000E-4   -3.990000E+2   -3.990000E+2   -6.319248E-2   -9.226258E-2   -1.407799E-4   -5.634555E-5   -1.407791E-4   -5.634776E-5   1.516371E-4   -1.581868E+2   -1.581859E+2   
3.349000E+3   2.028329E+1   2.028329E+1   -4.090000E+2   -4.090000E+2   9.000000E-4   -4.090000E+2   -4.090000E+2   -6.418702E-2   -9.108460E-2   -1.413062E-4   -5.770289E-5   -1.413053E-4   -5.770511E-5   1.526337E-4   -1.577872E+2   -1.577863E+2   
3.375796E+3   2.025860E+1   2.025860E+1   -4.190000E+2   -4.190000E+2   9.000000E-4   -4.190000E+2   -4.190000E+2   -6.459456E-2   -9.305831E-2   -1.436411E-4   -5.672089E-5   -1.436402E-4   -5.672315E-5   1.544345E-4   -1.584520E+2   -1.584511E+2   
3.402614E+3   2.025591E+1   2.025591E+1   -4.290000E+2   -4.290000E+2   9.000000E-4   -4.280000E+2   -4.280000E+2   -6.463385E-2   -9.617708E-2   -1.464591E-4   -5.478897E-5   -1.464582E-4   -5.479127E-5   1.563716E-4   -1.594896E+2   -1.594887E+2   
3.429400E+3   2.026431E+1   2.026431E+1   -4.390000E+2   -4.390000E+2   9.000000E-4   -4.380000E+2   -4.380000E+2   -6.528409E-2   -9.734911E-2   -1.483988E-4   -5.446435E-5   -1.483979E-4   -5.446668E-5   1.580777E-4   -1.598462E+2   -1.598453E+2   
3.456208E+3   2.025311E+1   2.025311E+1   -4.490000E+2   -4.490000E+2   9.000000E-4   -4.480000E+2   -4.480000E+2   -6.693113E-2   -9.856837E-2   -1.510642E-4   -5.477583E-5   -1.510633E-4   -5.477821E-5   1.606884E-4   -1.600694E+2   -1.600685E+2   
3.482995E+3   2.026309E+1   2.026309E+1   -4.590000E+2   -4.590000E+2   9.000000E-4   -4.580000E+2   -4.580000E+2   -6.862040E-2   -9.845961E-2   -1.528249E-4   -5.593615E-5   -1.528241E-4   -5.593855E-5   1.627400E-4   -1.598966E+2   -1.598957E+2   
3.509805E+3   2.027300E+1   2.027300E+1   -4.690000E+2   -4.690000E+2   9.000000E-4   -4.690000E+2   -4.690000E+2   -6.829969E-2   -1.021099E-1   -1.558994E-4   -5.342862E-5   -1.558986E-4   -5.343107E-5   1.648006E-4   -1.610828E+2   -1.610819E+2   
3.536617E+3   2.026409E+1   2.026409E+1   -4.790000E+2   -4.790000E+2   9.000000E-4   -4.780000E+2   -4.780000E+2   -6.937147E-2   -1.020892E-1   -1.572268E-4   -5.412581E-5   -1.572259E-4   -5.412828E-5   1.662825E-4   -1.610038E+2   -1.610029E+2   
3.563404E+3   2.028011E+1   2.028011E+1   -4.890000E+2   -4.890000E+2   9.000000E-4   -4.880000E+2   -4.880000E+2   -6.977840E-2   -1.014601E-1   -1.577308E-4   -5.475179E-5   -1.577300E-4   -5.475426E-5   1.669634E-4   -1.608570E+2   -1.608561E+2   
3.590215E+3   2.027041E+1   2.027041E+1   -4.990000E+2   -4.990000E+2   9.000000E-4   -4.980000E+2   -4.980000E+2   -7.114602E-2   -1.035735E-1   -1.608309E-4   -5.432430E-5   -1.608300E-4   -5.432683E-5   1.697577E-4   -1.613364E+2   -1.613355E+2   
3.617010E+3   2.028289E+1   2.028289E+1   -5.090000E+2   -5.090000E+2   9.000000E-4   -5.080000E+2   -5.080000E+2   -7.306182E-2   -1.033748E-1   -1.626857E-4   -5.569138E-5   -1.626849E-4   -5.569393E-5   1.719540E-4   -1.611026E+2   -1.611017E+2   
3.643802E+3   2.029019E+1   2.029019E+1   -5.190000E+2   -5.190000E+2   9.000000E-4   -5.180000E+2   -5.180000E+2   -7.271265E-2   -1.034872E-1   -1.631860E-4   -5.535446E-5   -1.631852E-4   -5.535703E-5   1.723189E-4   -1.612625E+2   -1.612616E+2   
3.670618E+3   2.029019E+1   2.029019E+1   -5.290000E+2   -5.290000E+2   9.000000E-4   -5.280000E+2   -5.280000E+2   -7.417536E-2   -1.068158E-1   -1.672068E-4   -5.423950E-5   -1.672059E-4   -5.424213E-5   1.757840E-4   -1.620277E+2   -1.620268E+2   
3.697425E+3   2.030490E+1   2.030490E+1   -5.390000E+2   -5.390000E+2   9.000000E-4   -5.380000E+2   -5.380000E+2   -7.405607E-2   -1.075797E-1   -1.683249E-4   -5.365348E-5   -1.683240E-4   -5.365612E-5   1.766691E-4   -1.623203E+2   -1.623194E+2   
3.724215E+3   2.029510E+1   2.029510E+1   -5.490000E+2   -5.490000E+2   9.000000E-4   -5.480000E+2   -5.480000E+2   -7.520371E-2   -1.096183E-1   -1.712196E-4   -5.312534E-5   -1.712187E-4   -5.312803E-5   1.792720E-4   -1.627621E+2   -1.627612E+2   
3.751004E+3   2.030499E+1   2.030499E+1   -5.590000E+2   -5.590000E+2   9.000000E-4   -5.580000E+2   -5.580000E+2   -7.650555E-2   -1.118050E-1   -1.743255E-4   -5.260863E-5   -1.743246E-4   -5.261137E-5   1.820907E-4   -1.632070E+2   -1.632061E+2   
3.777814E+3   2.029800E+1   2.029800E+1   -5.690000E+2   -5.690000E+2   9.000000E-4   -5.680000E+2   -5.680000E+2   -7.652687E-2   -1.116614E-1   -1.749031E-4   -5.267719E-5   -1.749023E-4   -5.267994E-5   1.826636E-4   -1.632388E+2   -1.632379E+2   
3.804620E+3   2.030529E+1   2.030529E+1   -5.790000E+2   -5.790000E+2   9.000000E-4   -5.790000E+2   -5.790000E+2   -7.782229E-2   -1.122358E-1   -1.769371E-4   -5.314906E-5   -1.769362E-4   -5.315184E-5   1.847473E-4   -1.632806E+2   -1.632797E+2   
3.831397E+3   2.029421E+1   2.029421E+1   -5.890000E+2   -5.890000E+2   9.000000E-4   -5.880000E+2   -5.880000E+2   -7.831331E-2   -1.118997E-1   -1.776392E-4   -5.365352E-5   -1.776384E-4   -5.365631E-5   1.855651E-4   -1.631938E+2   -1.631929E+2   
3.858208E+3   2.029711E+1   2.029711E+1   -5.990000E+2   -5.990000E+2   9.000000E-4   -5.980000E+2   -5.980000E+2   -7.921097E-2   -1.147453E-1   -1.809277E-4   -5.245988E-5   -1.809269E-4   -5.246273E-5   1.883796E-4   -1.638305E+2   -1.638296E+2   
3.885017E+3   2.028671E+1   2.028671E+1   -6.090000E+2   -6.090000E+2   9.000000E-4   -6.080000E+2   -6.080000E+2   -7.982660E-2   -1.138861E-1   -1.814149E-4   -5.336737E-5   -1.814141E-4   -5.337022E-5   1.891017E-4   -1.636075E+2   -1.636066E+2   
3.911820E+3   2.028701E+1   2.028701E+1   -6.190000E+2   -6.190000E+2   9.000000E-4   -6.190000E+2   -6.190000E+2   -8.007615E-2   -1.149275E-1   -1.830508E-4   -5.285256E-5   -1.830500E-4   -5.285544E-5   1.905282E-4   -1.638949E+2   -1.638940E+2   
3.938619E+3   2.028179E+1   2.028179E+1   -6.290000E+2   -6.290000E+2   9.000000E-4   -6.290000E+2   -6.290000E+2   -8.298207E-2   -1.160034E-1   -1.864899E-4   -5.409286E-5   -1.864890E-4   -5.409579E-5   1.941765E-4   -1.638248E+2   -1.638239E+2   
3.965420E+3   2.029110E+1   2.029110E+1   -6.390000E+2   -6.390000E+2   9.000000E-4   -6.380000E+2   -6.380000E+2   -8.217949E-2   -1.193231E-1   -1.888644E-4   -5.147489E-5   -1.888635E-4   -5.147786E-5   1.957534E-4   -1.647544E+2   -1.647535E+2   
3.992217E+3   2.028439E+1   2.028439E+1   -6.490000E+2   -6.490000E+2   9.000000E-4   -6.490000E+2   -6.490000E+2   -8.209676E-2   -1.192125E-1   -1.894593E-4   -5.145021E-5   -1.894585E-4   -5.145318E-5   1.963210E-4   -1.648070E+2   -1.648061E+2   
4.019028E+3   2.030499E+1   2.030499E+1   -6.600000E+2   -6.600000E+2   9.000000E-4   -6.590000E+2   -6.590000E+2   -8.321380E-2   -1.207003E-1   -1.919453E-4   -5.124201E-5   -1.919445E-4   -5.124502E-5   1.986674E-4   -1.650528E+2   -1.650519E+2   
4.045823E+3   2.029659E+1   2.029659E+1   -6.700000E+2   -6.700000E+2   9.000000E-4   -6.690000E+2   -6.690000E+2   -8.333034E-2   -1.199203E-1   -1.921415E-4   -5.176743E-5   -1.921407E-4   -5.177045E-5   1.989930E-4   -1.649212E+2   -1.649203E+2   
4.072608E+3   2.028500E+1   2.028500E+1   -6.790000E+2   -6.790000E+2   9.000000E-4   -6.790000E+2   -6.790000E+2   -8.426107E-2   -1.208469E-1   -1.941035E-4   -5.178168E-5   -1.941026E-4   -5.178473E-5   2.008917E-4   -1.650629E+2   -1.650620E+2   
4.099410E+3   2.030920E+1   2.030920E+1   -6.900000E+2   -6.900000E+2   9.000000E-4   -6.890000E+2   -6.890000E+2   -8.428194E-2   -1.216766E-1   -1.953652E-4   -5.124854E-5   -1.953644E-4   -5.125161E-5   2.019752E-4   -1.653013E+2   -1.653004E+2   
4.126209E+3   2.029650E+1   2.029650E+1   -6.990000E+2   -6.990000E+2   9.000000E-4   -6.990000E+2   -6.990000E+2   -8.526688E-2   -1.219740E-1   -1.969223E-4   -5.168778E-5   -1.969215E-4   -5.169087E-5   2.035928E-4   -1.652929E+2   -1.652920E+2   
4.153010E+3   2.029510E+1   2.029510E+1   -7.100000E+2   -7.100000E+2   9.000000E-4   -7.090000E+2   -7.090000E+2   -8.624314E-2   -1.243193E-1   -1.999136E-4   -5.085576E-5   -1.999128E-4   -5.085890E-5   2.062808E-4   -1.657273E+2   -1.657264E+2   
4.179802E+3   2.030529E+1   2.030529E+1   -7.200000E+2   -7.200000E+2   9.000000E-4   -7.190000E+2   -7.190000E+2   -8.684903E-2   -1.257794E-1   -2.020251E-4   -5.032353E-5   -2.020243E-4   -5.032670E-5   2.081985E-4   -1.660125E+2   -1.660116E+2   
4.206601E+3   2.030999E+1   2.030999E+1   -7.300000E+2   -7.300000E+2   9.000000E-4   -7.290000E+2   -7.290000E+2   -8.865852E-2   -1.251986E-1   -2.035375E-4   -5.185574E-5   -2.035367E-4   -5.185893E-5   2.100393E-4   -1.657067E+2   -1.657058E+2   
4.233397E+3   2.031521E+1   2.031521E+1   -7.400000E+2   -7.400000E+2   9.000000E-4   -7.390000E+2   -7.390000E+2   -8.967321E-2   -1.232502E-1   -2.035359E-4   -5.370261E-5   -2.035350E-4   -5.370580E-5   2.105014E-4   -1.652194E+2   -1.652185E+2   
4.260189E+3   2.031979E+1   2.031979E+1   -7.500000E+2   -7.500000E+2   9.000000E-4   -7.490000E+2   -7.490000E+2   -8.936942E-2   -1.272508E-1   -2.068021E-4   -5.099337E-5   -2.068013E-4   -5.099662E-5   2.129963E-4   -1.661483E+2   -1.661474E+2   
4.287022E+3   2.032171E+1   2.032171E+1   -7.590000E+2   -7.590000E+2   9.000000E-4   -7.590000E+2   -7.590000E+2   -8.777125E-2   -1.314443E-1   -2.093048E-4   -4.730097E-5   -2.093040E-4   -4.730426E-5   2.145830E-4   -1.672656E+2   -1.672647E+2   
4.313823E+3   2.032870E+1   2.032870E+1   -7.690000E+2   -7.690000E+2   9.000000E-4   -7.680000E+2   -7.680000E+2   -8.940812E-2   -1.295570E-1   -2.097120E-4   -4.952879E-5   -2.097112E-4   -4.953208E-5   2.154814E-4   -1.667117E+2   -1.667108E+2   
4.340625E+3   2.032510E+1   2.032510E+1   -7.790000E+2   -7.790000E+2   9.000000E-4   -7.790000E+2   -7.790000E+2   -9.052426E-2   -1.294112E-1   -2.111150E-4   -5.032600E-5   -2.111142E-4   -5.032932E-5   2.170305E-4   -1.665920E+2   -1.665911E+2   
4.367422E+3   2.032531E+1   2.032531E+1   -7.890000E+2   -7.890000E+2   9.000000E-4   -7.890000E+2   -7.890000E+2   -9.076585E-2   -1.311500E-1   -2.131694E-4   -4.937843E-5   -2.131686E-4   -4.938178E-5   2.188136E-4   -1.669581E+2   -1.669572E+2   
4.394222E+3   2.033749E+1   2.033749E+1   -7.990000E+2   -7.990000E+2   9.000000E-4   -7.990000E+2   -7.990000E+2   -9.298199E-2   -1.344083E-1   -2.176640E-4   -4.880976E-5   -2.176633E-4   -4.881318E-5   2.230696E-4   -1.673609E+2   -1.673600E+2   
4.421018E+3   2.032659E+1   2.032659E+1   -8.090000E+2   -8.090000E+2   9.000000E-4   -8.090000E+2   -8.090000E+2   -9.202109E-2   -1.349115E-1   -2.180142E-4   -4.782309E-5   -2.180135E-4   -4.782652E-5   2.231978E-4   -1.676277E+2   -1.676268E+2   
4.447819E+3   2.034231E+1   2.034231E+1   -8.190000E+2   -8.190000E+2   9.000000E-4   -8.190000E+2   -8.190000E+2   -9.451569E-2   -1.327361E-1   -2.188810E-4   -5.079797E-5   -2.188802E-4   -5.080140E-5   2.246983E-4   -1.669341E+2   -1.669332E+2   
4.474624E+3   2.033721E+1   2.033721E+1   -8.290000E+2   -8.290000E+2   9.000000E-4   -8.290000E+2   -8.290000E+2   -9.390037E-2   -1.360918E-1   -2.214772E-4   -4.827932E-5   -2.214765E-4   -4.828280E-5   2.266783E-4   -1.677026E+2   -1.677017E+2   
4.501421E+3   2.032711E+1   2.032711E+1   -8.390000E+2   -8.390000E+2   9.000000E-4   -8.390000E+2   -8.390000E+2   -9.524122E-2   -1.363308E-1   -2.232406E-4   -4.899217E-5   -2.232398E-4   -4.899568E-5   2.285532E-4   -1.676221E+2   -1.676212E+2   
4.528222E+3   2.033920E+1   2.033920E+1   -8.500000E+2   -8.500000E+2   9.000000E-4   -8.490000E+2   -8.490000E+2   -9.564923E-2   -1.354638E-1   -2.235780E-4   -4.976590E-5   -2.235772E-4   -4.976941E-5   2.290497E-4   -1.674512E+2   -1.674503E+2   
4.555025E+3   2.033691E+1   2.033691E+1   -8.590000E+2   -8.590000E+2   9.000000E-4   -8.590000E+2   -8.590000E+2   -9.563811E-2   -1.383340E-1   -2.262526E-4   -4.795045E-5   -2.262519E-4   -4.795400E-5   2.312780E-4   -1.680342E+2   -1.680333E+2   
4.581822E+3   2.033691E+1   2.033691E+1   -8.690000E+2   -8.690000E+2   9.000000E-4   -8.690000E+2   -8.690000E+2   -9.617744E-2   -1.379237E-1   -2.270025E-4   -4.852959E-5   -2.270018E-4   -4.853315E-5   2.321320E-4   -1.679327E+2   -1.679318E+2   
4.608618E+3   2.032580E+1   2.032580E+1   -8.790000E+2   -8.790000E+2   9.000000E-4   -8.790000E+2   -8.790000E+2   -9.655297E-2   -1.396346E-1   -2.291304E-4   -4.768862E-5   -2.291296E-4   -4.769222E-5   2.340404E-4   -1.682429E+2   -1.682420E+2   
4.635423E+3   2.033120E+1   2.033120E+1   -8.890000E+2   -8.890000E+2   9.000000E-4   -8.890000E+2   -8.890000E+2   -9.746911E-2   -1.400036E-1   -2.306900E-4   -4.803771E-5   -2.306893E-4   -4.804133E-5   2.356385E-4   -1.682371E+2   -1.682362E+2   
4.662222E+3   2.031552E+1   2.031552E+1   -8.990000E+2   -8.990000E+2   9.000000E-4   -8.990000E+2   -8.990000E+2   -9.917179E-2   -1.396441E-1   -2.322838E-4   -4.936194E-5   -2.322830E-4   -4.936559E-5   2.374707E-4   -1.680027E+2   -1.680018E+2   
4.689019E+3   2.032430E+1   2.032430E+1   -9.090000E+2   -9.090000E+2   9.000000E-4   -9.090000E+2   -9.090000E+2   -9.892011E-2   -1.408423E-1   -2.336154E-4   -4.841915E-5   -2.336146E-4   -4.842282E-5   2.385803E-4   -1.682907E+2   -1.682898E+2   
4.715816E+3   2.033029E+1   2.033029E+1   -9.190000E+2   -9.190000E+2   9.000000E-4   -9.190000E+2   -9.190000E+2   -9.913751E-2   -1.417010E-1   -2.350340E-4   -4.799929E-5   -2.350333E-4   -4.800298E-5   2.398852E-4   -1.684576E+2   -1.684567E+2   
4.742645E+3   2.032491E+1   2.032491E+1   -9.290000E+2   -9.290000E+2   9.000000E-4   -9.290000E+2   -9.290000E+2   -1.002868E-1   -1.421250E-1   -2.367944E-4   -4.847002E-5   -2.367936E-4   -4.847374E-5   2.417042E-4   -1.684318E+2   -1.684309E+2   
4.769435E+3   2.034149E+1   2.034149E+1   -9.390000E+2   -9.390000E+2   9.000000E-4   -9.390000E+2   -9.390000E+2   -9.915125E-2   -1.437842E-1   -2.378361E-4   -4.665243E-5   -2.378354E-4   -4.665616E-5   2.423685E-4   -1.689021E+2   -1.689012E+2   
4.796231E+3   2.034570E+1   2.034570E+1   -9.490000E+2   -9.490000E+2   9.000000E-4   -9.490000E+2   -9.490000E+2   -9.942925E-2   -1.454951E-1   -2.398962E-4   -4.574638E-5   -2.398955E-4   -4.575014E-5   2.442190E-4   -1.692038E+2   -1.692029E+2   
4.823028E+3   2.035671E+1   2.035671E+1   -9.590000E+2   -9.590000E+2   9.000000E-4   -9.580000E+2   -9.580000E+2   -1.024034E-1   -1.455277E-1   -2.425826E-4   -4.768037E-5   -2.425819E-4   -4.768418E-5   2.472241E-4   -1.688801E+2   -1.688792E+2   
4.849825E+3   2.035650E+1   2.035650E+1   -9.690000E+2   -9.690000E+2   9.000000E-4   -9.690000E+2   -9.690000E+2   -1.028293E-1   -1.427200E-1   -2.416341E-4   -4.966173E-5   -2.416333E-4   -4.966552E-5   2.466846E-4   -1.683860E+2   -1.683851E+2   
4.876625E+3   2.035470E+1   2.035470E+1   -9.790000E+2   -9.790000E+2   9.000000E-4   -9.790000E+2   -9.790000E+2   -1.017368E-1   -1.497601E-1   -2.464899E-4   -4.454785E-5   -2.464892E-4   -4.455172E-5   2.504831E-4   -1.697556E+2   -1.697547E+2   
4.903425E+3   2.037039E+1   2.037039E+1   -9.890000E+2   -9.890000E+2   9.000000E-4   -9.890000E+2   -9.890000E+2   -1.048954E-1   -1.463100E-1   -2.469216E-4   -4.875361E-5   -2.469208E-4   -4.875749E-5   2.516887E-4   -1.688309E+2   -1.688300E+2   
4.930224E+3   2.037020E+1   2.037020E+1   -9.990000E+2   -9.990000E+2   9.000000E-4   -9.980000E+2   -9.980000E+2   -1.008001E-1   -1.500144E-1   -2.472792E-4   -4.370026E-5   -2.472786E-4   -4.370414E-5   2.511110E-4   -1.699779E+2   -1.699770E+2   
4.957142E+3   2.036730E+1   2.036730E+1   -1.009000E+3   -1.009000E+3   9.000000E-4   -1.008000E+3   -1.008000E+3   -1.027911E-1   -1.516958E-1   -2.505086E-4   -4.395567E-5   -2.505079E-4   -4.395961E-5   2.543357E-4   -1.700479E+2   -1.700470E+2   
4.984097E+3   2.038040E+1   2.038040E+1   -1.019000E+3   -1.019000E+3   9.000000E-4   -1.019000E+3   -1.019000E+3   -1.037618E-1   -1.540705E-1   -2.535831E-4   -4.309837E-5   -2.535824E-4   -4.310235E-5   2.572195E-4   -1.703543E+2   -1.703534E+2   
5.011065E+3   2.037881E+1   2.037881E+1   -1.029000E+3   -1.029000E+3   9.000000E-4   -1.028000E+3   -1.028000E+3   -1.046300E-1   -1.508354E-1   -2.525085E-4   -4.564605E-5   -2.525078E-4   -4.565002E-5   2.566010E-4   -1.697533E+2   -1.697524E+2   
5.038012E+3   2.038461E+1   2.038461E+1   -1.039000E+3   -1.039000E+3   9.000000E-4   -1.038000E+3   -1.038000E+3   -1.056537E-1   -1.507561E-1   -2.538276E-4   -4.634386E-5   -2.538269E-4   -4.634785E-5   2.580237E-4   -1.696529E+2   -1.696520E+2   
5.064923E+3   2.039141E+1   2.039141E+1   -1.049000E+3   -1.049000E+3   9.000000E-4   -1.049000E+3   -1.049000E+3   -1.074193E-1   -1.505793E-1   -2.556599E-4   -4.759375E-5   -2.556591E-4   -4.759777E-5   2.600522E-4   -1.694545E+2   -1.694536E+2   
5.091866E+3   2.038070E+1   2.038070E+1   -1.059000E+3   -1.059000E+3   9.000000E-4   -1.059000E+3   -1.059000E+3   -1.060972E-1   -1.522661E-1   -2.565915E-4   -4.563465E-5   -2.565908E-4   -4.563868E-5   2.606180E-4   -1.699154E+2   -1.699145E+2   
5.118778E+3   2.038131E+1   2.038131E+1   -1.069000E+3   -1.069000E+3   9.000000E-4   -1.068000E+3   -1.068000E+3   -1.070597E-1   -1.519414E-1   -2.576292E-4   -4.644677E-5   -2.576285E-4   -4.645082E-5   2.617826E-4   -1.697802E+2   -1.697793E+2   
5.145726E+3   2.037869E+1   2.037869E+1   -1.079000E+3   -1.079000E+3   9.000000E-4   -1.078000E+3   -1.078000E+3   -1.080032E-1   -1.523170E-1   -2.592125E-4   -4.681005E-5   -2.592118E-4   -4.681412E-5   2.634052E-4   -1.697635E+2   -1.697626E+2   
5.172666E+3   2.037029E+1   2.037029E+1   -1.089000E+3   -1.089000E+3   9.000000E-4   -1.088000E+3   -1.088000E+3   -1.068385E-1   -1.535385E-1   -2.599263E-4   -4.524347E-5   -2.599256E-4   -4.524755E-5   2.638345E-4   -1.701259E+2   -1.701250E+2   
5.199592E+3   2.037121E+1   2.037121E+1   -1.099000E+3   -1.099000E+3   9.000000E-4   -1.098000E+3   -1.098000E+3   -1.067199E-1   -1.548321E-1   -2.614174E-4   -4.433055E-5   -2.614167E-4   -4.433466E-5   2.651495E-4   -1.703755E+2   -1.703746E+2   
5.226533E+3   2.037390E+1   2.037390E+1   -1.109000E+3   -1.109000E+3   9.000000E-4   -1.109000E+3   -1.109000E+3   -1.090986E-1   -1.545553E-1   -2.636053E-4   -4.605147E-5   -2.636046E-4   -4.605561E-5   2.675976E-4   -1.700905E+2   -1.700896E+2   
5.253453E+3   2.036959E+1   2.036959E+1   -1.119000E+3   -1.119000E+3   9.000000E-4   -1.118000E+3   -1.118000E+3   -1.091337E-1   -1.552037E-1   -2.646830E-4   -4.564325E-5   -2.646823E-4   -4.564741E-5   2.685897E-4   -1.702159E+2   -1.702150E+2   
5.280409E+3   2.035540E+1   2.035540E+1   -1.129000E+3   -1.129000E+3   9.000000E-4   -1.129000E+3   -1.129000E+3   -1.088332E-1   -1.560750E-1   -2.658172E-4   -4.486653E-5   -2.658165E-4   -4.487071E-5   2.695771E-4   -1.704195E+2   -1.704186E+2   
5.307320E+3   2.036620E+1   2.036620E+1   -1.139000E+3   -1.139000E+3   9.000000E-4   -1.139000E+3   -1.139000E+3   -1.095831E-1   -1.573672E-1   -2.679107E-4   -4.453413E-5   -2.679100E-4   -4.453834E-5   2.715868E-4   -1.705622E+2   -1.705613E+2   
5.334293E+3   2.036379E+1   2.036379E+1   -1.149000E+3   -1.149000E+3   9.000000E-4   -1.148000E+3   -1.148000E+3   -1.100360E-1   -1.565326E-1   -2.682358E-4   -4.532122E-5   -2.682351E-4   -4.532543E-5   2.720376E-4   -1.704099E+2   -1.704090E+2   
5.361332E+3   2.036321E+1   2.036321E+1   -1.159000E+3   -1.159000E+3   9.000000E-4   -1.158000E+3   -1.158000E+3   -1.101817E-1   -1.587513E-1   -2.705610E-4   -4.401304E-5   -2.705603E-4   -4.401729E-5   2.741175E-4   -1.707604E+2   -1.707595E+2   
5.388276E+3   2.036031E+1   2.036031E+1   -1.169000E+3   -1.169000E+3   9.000000E-4   -1.168000E+3   -1.168000E+3   -1.111771E-1   -1.593432E-1   -2.723325E-4   -4.427733E-5   -2.723319E-4   -4.428161E-5   2.759085E-4   -1.707653E+2   -1.707644E+2   
5.415323E+3   2.036208E+1   2.036208E+1   -1.179000E+3   -1.179000E+3   9.000000E-4   -1.178000E+3   -1.178000E+3   -1.109760E-1   -1.590433E-1   -2.726458E-4   -4.429402E-5   -2.726451E-4   -4.429830E-5   2.762203E-4   -1.707723E+2   -1.707714E+2   
5.442320E+3   2.035671E+1   2.035671E+1   -1.189000E+3   -1.189000E+3   9.000000E-4   -1.188000E+3   -1.188000E+3   -1.126065E-1   -1.600961E-1   -2.751825E-4   -4.469733E-5   -2.751818E-4   -4.470165E-5   2.787889E-4   -1.707741E+2   -1.707732E+2   
5.469322E+3   2.036599E+1   2.036599E+1   -1.199000E+3   -1.199000E+3   9.000000E-4   -1.198000E+3   -1.198000E+3   -1.121525E-1   -1.607427E-1   -2.759856E-4   -4.396040E-5   -2.759849E-4   -4.396473E-5   2.794648E-4   -1.709497E+2   -1.709488E+2   
5.496268E+3   2.036770E+1   2.036770E+1   -1.209000E+3   -1.209000E+3   9.000000E-4   -1.209000E+3   -1.209000E+3   -1.141319E-1   -1.610280E-1   -2.782915E-4   -4.506743E-5   -2.782908E-4   -4.507180E-5   2.819171E-4   -1.708012E+2   -1.708003E+2   
5.523222E+3   2.036700E+1   2.036700E+1   -1.219000E+3   -1.219000E+3   9.000000E-4   -1.218000E+3   -1.218000E+3   -1.133359E-1   -1.625043E-1   -2.793741E-4   -4.359297E-5   -2.793735E-4   -4.359735E-5   2.827548E-4   -1.711312E+2   -1.711303E+2   
5.550169E+3   2.036340E+1   2.036340E+1   -1.229000E+3   -1.229000E+3   9.000000E-4   -1.229000E+3   -1.229000E+3   -1.124669E-1   -1.628626E-1   -2.797526E-4   -4.275375E-5   -2.797519E-4   -4.275814E-5   2.830007E-4   -1.713109E+2   -1.713100E+2   
5.577188E+3   2.037911E+1   2.037911E+1   -1.239000E+3   -1.239000E+3   9.000000E-4   -1.238000E+3   -1.238000E+3   -1.139068E-1   -1.638384E-1   -2.820365E-4   -4.308082E-5   -2.820358E-4   -4.308525E-5   2.853078E-4   -1.713152E+2   -1.713143E+2   
5.604167E+3   2.037969E+1   2.037969E+1   -1.249000E+3   -1.249000E+3   9.000000E-4   -1.248000E+3   -1.248000E+3   -1.139557E-1   -1.618512E-1   -2.813367E-4   -4.430710E-5   -2.813360E-4   -4.431152E-5   2.848042E-4   -1.710501E+2   -1.710492E+2   
5.631072E+3   2.040679E+1   2.040679E+1   -1.259000E+3   -1.259000E+3   9.000000E-4   -1.258000E+3   -1.258000E+3   -1.145562E-1   -1.635686E-1   -2.836254E-4   -4.361230E-5   -2.836247E-4   -4.361676E-5   2.869589E-4   -1.712583E+2   -1.712574E+2   
5.657991E+3   2.040621E+1   2.040621E+1   -1.269000E+3   -1.269000E+3   9.000000E-4   -1.268000E+3   -1.268000E+3   -1.133768E-1   -1.652196E-1   -2.846310E-4   -4.177047E-5   -2.846303E-4   -4.177494E-5   2.876796E-4   -1.716513E+2   -1.716504E+2   
5.684992E+3   2.040759E+1   2.040759E+1   -1.278000E+3   -1.278000E+3   9.000000E-4   -1.278000E+3   -1.278000E+3   -1.159932E-1   -1.643684E-1   -2.865137E-4   -4.400837E-5   -2.865130E-4   -4.401287E-5   2.898738E-4   -1.712676E+2   -1.712667E+2   
5.712005E+3   2.042489E+1   2.042489E+1   -1.289000E+3   -1.289000E+3   9.000000E-4   -1.288000E+3   -1.288000E+3   -1.154423E-1   -1.650353E-1   -2.872637E-4   -4.319427E-5   -2.872630E-4   -4.319879E-5   2.904930E-4   -1.714488E+2   -1.714479E+2   
5.738951E+3   2.041781E+1   2.041781E+1   -1.299000E+3   -1.299000E+3   9.000000E-4   -1.298000E+3   -1.298000E+3   -1.162545E-1   -1.660039E-1   -2.891729E-4   -4.310341E-5   -2.891722E-4   -4.310795E-5   2.923677E-4   -1.715221E+2   -1.715212E+2   
5.765877E+3   2.040640E+1   2.040640E+1   -1.309000E+3   -1.309000E+3   9.000000E-4   -1.308000E+3   -1.308000E+3   -1.171806E-1   -1.679693E-1   -2.918622E-4   -4.247268E-5   -2.918615E-4   -4.247727E-5   2.949364E-4   -1.717203E+2   -1.717194E+2   
5.792816E+3   2.041360E+1   2.041360E+1   -1.319000E+3   -1.319000E+3   9.000000E-4   -1.318000E+3   -1.318000E+3   -1.161699E-1   -1.674763E-1   -2.914771E-4   -4.206840E-5   -2.914765E-4   -4.207298E-5   2.944973E-4   -1.717873E+2   -1.717864E+2   
5.819744E+3   2.041241E+1   2.041241E+1   -1.329000E+3   -1.329000E+3   9.000000E-4   -1.328000E+3   -1.328000E+3   -1.174411E-1   -1.684579E-1   -2.937143E-4   -4.227589E-5   -2.937137E-4   -4.228050E-5   2.967412E-4   -1.718094E+2   -1.718085E+2   
5.846691E+3   2.040688E+1   2.040688E+1   -1.339000E+3   -1.339000E+3   9.000000E-4   -1.338000E+3   -1.338000E+3   -1.185539E-1   -1.692200E-1   -2.956871E-4   -4.251325E-5   -2.956864E-4   -4.251790E-5   2.987277E-4   -1.718182E+2   -1.718173E+2   
5.873620E+3   2.040991E+1   2.040991E+1   -1.349000E+3   -1.349000E+3   9.000000E-4   -1.348000E+3   -1.348000E+3   -1.168337E-1   -1.698167E-1   -2.955755E-4   -4.096210E-5   -2.955748E-4   -4.096674E-5   2.984003E-4   -1.721100E+2   -1.721091E+2   
5.900562E+3   2.041351E+1   2.041351E+1   -1.359000E+3   -1.359000E+3   9.000000E-4   -1.358000E+3   -1.358000E+3   -1.198010E-1   -1.688414E-1   -2.976147E-4   -4.351084E-5   -2.976140E-4   -4.351552E-5   3.007785E-4   -1.716824E+2   -1.716815E+2   
5.927516E+3   2.040771E+1   2.040771E+1   -1.369000E+3   -1.369000E+3   9.000000E-4   -1.368000E+3   -1.368000E+3   -1.195396E-1   -1.696669E-1   -2.986774E-4   -4.279189E-5   -2.986767E-4   -4.279658E-5   3.017273E-4   -1.718466E+2   -1.718457E+2   
5.954537E+3   2.040209E+1   2.040209E+1   -1.379000E+3   -1.379000E+3   9.000000E-4   -1.378000E+3   -1.378000E+3   -1.199942E-1   -1.696089E-1   -2.996162E-4   -4.309683E-5   -2.996155E-4   -4.310153E-5   3.026998E-4   -1.718147E+2   -1.718138E+2   
5.981527E+3   2.039019E+1   2.039019E+1   -1.389000E+3   -1.389000E+3   9.000000E-4   -1.388000E+3   -1.388000E+3   -1.195052E-1   -1.717314E-1   -3.014329E-4   -4.142444E-5   -3.014323E-4   -4.142918E-5   3.042660E-4   -1.721751E+2   -1.721742E+2   
6.008432E+3   2.039660E+1   2.039660E+1   -1.399000E+3   -1.399000E+3   9.000000E-4   -1.398000E+3   -1.398000E+3   -1.200794E-1   -1.712043E-1   -3.021249E-4   -4.209905E-5   -3.021242E-4   -4.210380E-5   3.050439E-4   -1.720673E+2   -1.720664E+2   
6.035373E+3   2.039309E+1   2.039309E+1   -1.409000E+3   -1.409000E+3   9.000000E-4   -1.408000E+3   -1.408000E+3   -1.207589E-1   -1.722478E-1   -3.039945E-4   -4.187340E-5   -3.039938E-4   -4.187818E-5   3.068648E-4   -1.721572E+2   -1.721563E+2   
6.062320E+3   2.038879E+1   2.038879E+1   -1.419000E+3   -1.419000E+3   9.000000E-4   -1.418000E+3   -1.418000E+3   -1.207811E-1   -1.739541E-1   -3.058737E-4   -4.079946E-5   -3.058730E-4   -4.080426E-5   3.085827E-4   -1.724024E+2   -1.724015E+2   
6.089328E+3   2.039419E+1   2.039419E+1   -1.429000E+3   -1.429000E+3   9.000000E-4   -1.428000E+3   -1.428000E+3   -1.211347E-1   -1.742794E-1   -3.070119E-4   -4.080010E-5   -3.070112E-4   -4.080493E-5   3.097110E-4   -1.724301E+2   -1.724292E+2   
6.116289E+3   2.039471E+1   2.039471E+1   -1.439000E+3   -1.439000E+3   9.000000E-4   -1.438000E+3   -1.438000E+3   -1.220878E-1   -1.758986E-1   -3.094764E-4   -4.040129E-5   -3.094758E-4   -4.040616E-5   3.121024E-4   -1.725623E+2   -1.725614E+2   
6.143233E+3   2.039239E+1   2.039239E+1   -1.449000E+3   -1.449000E+3   9.000000E-4   -1.448000E+3   -1.448000E+3   -1.208845E-1   -1.744211E-1   -3.082653E-4   -4.047683E-5   -3.082646E-4   -4.048168E-5   3.109113E-4   -1.725196E+2   -1.725187E+2   
6.170176E+3   2.038000E+1   2.038000E+1   -1.459000E+3   -1.459000E+3   9.000000E-4   -1.458000E+3   -1.458000E+3   -1.229368E-1   -1.747672E-1   -3.105981E-4   -4.159835E-5   -3.105975E-4   -4.160323E-5   3.133714E-4   -1.723718E+2   -1.723709E+2   
6.197067E+3   2.039419E+1   2.039419E+1   -1.469000E+3   -1.469000E+3   9.000000E-4   -1.468000E+3   -1.468000E+3   -1.236972E-1   -1.754473E-1   -3.122684E-4   -4.165123E-5   -3.122677E-4   -4.165614E-5   3.150339E-4   -1.724026E+2   -1.724017E+2   
6.224027E+3   2.039099E+1   2.039099E+1   -1.479000E+3   -1.479000E+3   9.000000E-4   -1.478000E+3   -1.478000E+3   -1.216177E-1   -1.766800E-1   -3.123545E-4   -3.946718E-5   -3.123538E-4   -3.947208E-5   3.148380E-4   -1.727986E+2   -1.727977E+2   
6.250959E+3   2.040911E+1   2.040911E+1   -1.489000E+3   -1.489000E+3   9.000000E-4   -1.488000E+3   -1.488000E+3   -1.223079E-1   -1.802051E-1   -3.159768E-4   -3.771522E-5   -3.159762E-4   -3.772018E-5   3.182197E-4   -1.731933E+2   -1.731924E+2   
6.277929E+3   2.041580E+1   2.041580E+1   -1.498000E+3   -1.498000E+3   9.000000E-4   -1.498000E+3   -1.498000E+3   -1.216234E-1   -1.794100E-1   -3.156059E-4   -3.771528E-5   -3.156054E-4   -3.772024E-5   3.178515E-4   -1.731854E+2   -1.731845E+2   
6.304966E+3   2.041729E+1   2.041729E+1   -1.509000E+3   -1.509000E+3   9.000000E-4   -1.508000E+3   -1.508000E+3   -1.234210E-1   -1.893997E-1   -3.245437E-4   -3.270767E-5   -3.245432E-4   -3.271277E-5   3.261877E-4   -1.742451E+2   -1.742442E+2   
6.332672E+3   2.043209E+1   2.043209E+1   -1.518000E+3   -1.518000E+3   9.000000E-4   -1.518000E+3   -1.518000E+3   -1.260374E-1   -1.803567E-1   -3.206655E-4   -4.000761E-5   -3.206649E-4   -4.001265E-5   3.231517E-4   -1.728883E+2   -1.728874E+2   
6.359645E+3   2.043301E+1   2.043301E+1   -1.529000E+3   -1.529000E+3   9.000000E-4   -1.528000E+3   -1.528000E+3   -1.275955E-1   -1.753310E-1   -3.188773E-4   -4.411873E-5   -3.188766E-4   -4.412374E-5   3.219149E-4   -1.721228E+2   -1.721219E+2   
6.387080E+3   2.043249E+1   2.043249E+1   -1.539000E+3   -1.539000E+3   9.000000E-4   -1.538000E+3   -1.538000E+3   -1.241351E-1   -1.787420E-1   -3.195360E-4   -3.966695E-5   -3.195354E-4   -3.967197E-5   3.219887E-4   -1.729235E+2   -1.729226E+2   
6.414050E+3   2.043780E+1   2.043780E+1   -1.548000E+3   -1.548000E+3   9.000000E-4   -1.548000E+3   -1.548000E+3   -1.247205E-1   -1.794009E-1   -3.210699E-4   -3.961617E-5   -3.210693E-4   -3.962121E-5   3.235047E-4   -1.729659E+2   -1.729650E+2   
6.441728E+3   2.042590E+1   2.042590E+1   -1.559000E+3   -1.559000E+3   9.000000E-4   -1.557000E+3   -1.557000E+3   -1.261118E-1   -1.794442E-1   -3.226642E-4   -4.048707E-5   -3.226636E-4   -4.049214E-5   3.251944E-4   -1.728481E+2   -1.728472E+2   
6.468702E+3   2.041189E+1   2.041189E+1   -1.568000E+3   -1.568000E+3   9.000000E-4   -1.568000E+3   -1.568000E+3   -1.244075E-1   -1.791218E-1   -3.219836E-4   -3.951097E-5   -3.219830E-4   -3.951603E-5   3.243988E-4   -1.730041E+2   -1.730032E+2   
6.496368E+3   2.042281E+1   2.042281E+1   -1.579000E+3   -1.579000E+3   9.000000E-4   -1.578000E+3   -1.578000E+3   -1.397853E-1   -1.778568E-1   -3.324403E-4   -5.052195E-5   -3.324395E-4   -5.052717E-5   3.362574E-4   -1.713587E+2   -1.713578E+2   
6.523395E+3   2.044070E+1   2.044070E+1   -1.589000E+3   -1.589000E+3   9.000000E-4   -1.588000E+3   -1.588000E+3   -1.247653E-1   -1.953009E-1   -3.349379E-4   -2.968339E-5   -3.349374E-4   -2.968865E-5   3.362506E-4   -1.749355E+2   -1.749346E+2   
6.550438E+3   2.043279E+1   2.043279E+1   -1.598000E+3   -1.598000E+3   9.000000E-4   -1.597000E+3   -1.597000E+3   -1.275856E-1   -1.839598E-1   -3.295187E-4   -3.854293E-5   -3.295181E-4   -3.854811E-5   3.317652E-4   -1.733286E+2   -1.733277E+2   
6.577831E+3   2.043051E+1   2.043051E+1   -1.609000E+3   -1.609000E+3   9.000000E-4   -1.608000E+3   -1.608000E+3   -1.240865E-1   -1.783634E-1   -3.238824E-4   -3.962790E-5   -3.238818E-4   -3.963299E-5   3.262977E-4   -1.730244E+2   -1.730235E+2   
6.604873E+3   2.042870E+1   2.042870E+1   -1.619000E+3   -1.619000E+3   9.000000E-4   -1.618000E+3   -1.618000E+3   -1.249754E-1   -1.832439E-1   -3.285959E-4   -3.717102E-5   -3.285954E-4   -3.717619E-5   3.306917E-4   -1.735461E+2   -1.735452E+2   
6.632598E+3   2.043710E+1   2.043710E+1   -1.629000E+3   -1.629000E+3   9.000000E-4   -1.628000E+3   -1.628000E+3   -1.315601E-1   -2.067011E-1   -3.503304E-4   -2.703630E-5   -3.503300E-4   -2.704181E-5   3.513721E-4   -1.755870E+2   -1.755861E+2   
6.659514E+3   2.043041E+1   2.043041E+1   -1.638000E+3   -1.638000E+3   9.000000E-4   -1.637000E+3   -1.637000E+3   -1.282654E-1   -1.865873E-1   -3.344939E-4   -3.723549E-5   -3.344933E-4   -3.724075E-5   3.365600E-4   -1.736480E+2   -1.736471E+2   
6.686960E+3   2.043719E+1   2.043719E+1   -1.648000E+3   -1.648000E+3   9.000000E-4   -1.648000E+3   -1.648000E+3   -1.282051E-1   -1.833401E-1   -3.328985E-4   -3.916402E-5   -3.328979E-4   -3.916925E-5   3.351943E-4   -1.732902E+2   -1.732893E+2   
6.713896E+3   2.041931E+1   2.041931E+1   -1.658000E+3   -1.658000E+3   9.000000E-4   -1.658000E+3   -1.658000E+3   -1.301247E-1   -1.901858E-1   -3.397100E-4   -3.618066E-5   -3.397094E-4   -3.618599E-5   3.416313E-4   -1.739207E+2   -1.739198E+2   
6.740857E+3   2.041491E+1   2.041491E+1   -1.668000E+3   -1.668000E+3   9.000000E-4   -1.668000E+3   -1.668000E+3   -1.328519E-1   -1.896857E-1   -3.419166E-4   -3.827550E-5   -3.419160E-4   -3.828087E-5   3.440523E-4   -1.736127E+2   -1.736118E+2   
6.769095E+3   2.042260E+1   2.042260E+1   -1.678000E+3   -1.678000E+3   9.000000E-4   -1.677000E+3   -1.677000E+3   -1.324398E-1   -1.890296E-1   -3.417663E-4   -3.837497E-5   -3.417657E-4   -3.838034E-5   3.439140E-4   -1.735934E+2   -1.735925E+2   
6.797032E+3   2.042529E+1   2.042529E+1   -1.689000E+3   -1.689000E+3   9.000000E-4   -1.688000E+3   -1.688000E+3   -1.320780E-1   -1.899836E-1   -3.429160E-4   -3.750612E-5   -3.429155E-4   -3.751151E-5   3.449610E-4   -1.737581E+2   -1.737572E+2   
6.824056E+3   2.042669E+1   2.042669E+1   -1.698000E+3   -1.698000E+3   9.000000E-4   -1.698000E+3   -1.698000E+3   -1.331398E-1   -1.902996E-1   -3.445397E-4   -3.798525E-5   -3.445391E-4   -3.799067E-5   3.466273E-4   -1.737086E+2   -1.737077E+2   
6.850987E+3   2.040869E+1   2.040869E+1   -1.708000E+3   -1.708000E+3   9.000000E-4   -1.708000E+3   -1.708000E+3   -1.350271E-1   -1.934621E-1   -3.487386E-4   -3.725626E-5   -3.487380E-4   -3.726173E-5   3.507230E-4   -1.739021E+2   -1.739012E+2   
6.879173E+3   2.041860E+1   2.041860E+1   -1.718000E+3   -1.718000E+3   9.000000E-4   -1.718000E+3   -1.718000E+3   -1.352644E-1   -1.938212E-1   -3.498197E-4   -3.715834E-5   -3.498191E-4   -3.716383E-5   3.517876E-4   -1.739367E+2   -1.739358E+2   
6.907421E+3   2.041921E+1   2.041921E+1   -1.728000E+3   -1.728000E+3   9.000000E-4   -1.727000E+3   -1.727000E+3   -1.363456E-1   -1.940106E-1   -3.513013E-4   -3.773203E-5   -3.513007E-4   -3.773755E-5   3.533218E-4   -1.738696E+2   -1.738687E+2   
6.934427E+3   2.042761E+1   2.042761E+1   -1.738000E+3   -1.738000E+3   9.000000E-4   -1.737000E+3   -1.737000E+3   -1.337351E-1   -1.981305E-1   -3.530490E-4   -3.340945E-5   -3.530485E-4   -3.341499E-5   3.546263E-4   -1.745941E+2   -1.745932E+2   
6.961380E+3   2.041311E+1   2.041311E+1   -1.748000E+3   -1.748000E+3   9.000000E-4   -1.748000E+3   -1.748000E+3   -1.366815E-1   -1.948467E-1   -3.535166E-4   -3.736739E-5   -3.535160E-4   -3.737295E-5   3.554860E-4   -1.739661E+2   -1.739652E+2   
6.989621E+3   2.040991E+1   2.040991E+1   -1.758000E+3   -1.758000E+3   9.000000E-4   -1.757000E+3   -1.757000E+3   -1.396932E-1   -1.977633E-1   -3.582573E-4   -3.754423E-5   -3.582567E-4   -3.754986E-5   3.602191E-4   -1.740174E+2   -1.740165E+2   
7.016622E+3   2.043621E+1   2.043621E+1   -1.768000E+3   -1.768000E+3   9.000000E-4   -1.768000E+3   -1.768000E+3   -1.332442E-1   -1.999733E-1   -3.560617E-4   -3.183657E-5   -3.560612E-4   -3.184216E-5   3.574822E-4   -1.748906E+2   -1.748897E+2   
7.043626E+3   2.043099E+1   2.043099E+1   -1.778000E+3   -1.778000E+3   9.000000E-4   -1.777000E+3   -1.777000E+3   -1.352034E-1   -2.110569E-1   -3.658147E-4   -2.626426E-5   -3.658143E-4   -2.627001E-5   3.667564E-4   -1.758934E+2   -1.758925E+2   
7.071862E+3   2.043411E+1   2.043411E+1   -1.788000E+3   -1.788000E+3   9.000000E-4   -1.787000E+3   -1.787000E+3   -1.373343E-1   -1.993504E-1   -3.597261E-4   -3.488607E-5   -3.597255E-4   -3.489172E-5   3.614137E-4   -1.744608E+2   -1.744599E+2   
7.100140E+3   2.043450E+1   2.043450E+1   -1.798000E+3   -1.798000E+3   9.000000E-4   -1.797000E+3   -1.797000E+3   -1.374792E-1   -1.980545E-1   -3.595792E-4   -3.574917E-5   -3.595786E-4   -3.575482E-5   3.613519E-4   -1.743223E+2   -1.743214E+2   
7.127130E+3   2.043530E+1   2.043530E+1   -1.808000E+3   -1.808000E+3   9.000000E-4   -1.807000E+3   -1.807000E+3   -1.379850E-1   -1.985256E-1   -3.609256E-4   -3.576127E-5   -3.609250E-4   -3.576694E-5   3.626929E-4   -1.743415E+2   -1.743406E+2   
7.154071E+3   2.043621E+1   2.043621E+1   -1.818000E+3   -1.818000E+3   9.000000E-4   -1.817000E+3   -1.817000E+3   -1.371303E-1   -2.008732E-1   -3.626466E-4   -3.370579E-5   -3.626461E-4   -3.371149E-5   3.642096E-4   -1.746900E+2   -1.746891E+2   
7.181469E+3   2.045669E+1   2.045669E+1   -1.828000E+3   -1.828000E+3   9.000000E-4   -1.827000E+3   -1.827000E+3   -1.387117E-1   -1.989396E-1   -3.630491E-4   -3.592177E-5   -3.630485E-4   -3.592747E-5   3.648219E-4   -1.743493E+2   -1.743484E+2   
7.209723E+3   2.044891E+1   2.044891E+1   -1.838000E+3   -1.838000E+3   9.000000E-4   -1.837000E+3   -1.837000E+3   -1.393545E-1   -1.990169E-1   -3.642138E-4   -3.626859E-5   -3.642132E-4   -3.627432E-5   3.660151E-4   -1.743132E+2   -1.743123E+2   
7.236725E+3   2.044659E+1   2.044659E+1   -1.848000E+3   -1.848000E+3   9.000000E-4   -1.847000E+3   -1.847000E+3   -1.376073E-1   -1.985254E-1   -3.633182E-4   -3.537184E-5   -3.633177E-4   -3.537755E-5   3.650360E-4   -1.744393E+2   -1.744384E+2   
7.263721E+3   2.044351E+1   2.044351E+1   -1.858000E+3   -1.858000E+3   9.000000E-4   -1.857000E+3   -1.857000E+3   -1.381098E-1   -1.999996E-1   -3.653678E-4   -3.476184E-5   -3.653672E-4   -3.476758E-5   3.670177E-4   -1.745651E+2   -1.745642E+2   
7.291210E+3   2.043389E+1   2.043389E+1   -1.868000E+3   -1.868000E+3   9.000000E-4   -1.867000E+3   -1.867000E+3   -1.384407E-1   -2.014693E-1   -3.672950E-4   -3.404015E-5   -3.672945E-4   -3.404592E-5   3.688690E-4   -1.747051E+2   -1.747042E+2   
7.319434E+3   2.042471E+1   2.042471E+1   -1.878000E+3   -1.878000E+3   9.000000E-4   -1.877000E+3   -1.877000E+3   -1.386794E-1   -2.010670E-1   -3.678416E-4   -3.441375E-5   -3.678411E-4   -3.441953E-5   3.694479E-4   -1.746552E+2   -1.746543E+2   
7.346427E+3   2.042840E+1   2.042840E+1   -1.888000E+3   -1.888000E+3   9.000000E-4   -1.887000E+3   -1.887000E+3   -1.396116E-1   -2.018510E-1   -3.697044E-4   -3.451709E-5   -3.697039E-4   -3.452290E-5   3.713122E-4   -1.746661E+2   -1.746652E+2   
7.373410E+3   2.043481E+1   2.043481E+1   -1.898000E+3   -1.898000E+3   9.000000E-4   -1.897000E+3   -1.897000E+3   -1.406007E-1   -1.989966E-1   -3.690478E-4   -3.690674E-5   -3.690472E-4   -3.691254E-5   3.708886E-4   -1.742891E+2   -1.742882E+2   
7.401586E+3   2.042849E+1   2.042849E+1   -1.908000E+3   -1.908000E+3   9.000000E-4   -1.907000E+3   -1.907000E+3   -1.368965E-1   -2.023012E-1   -3.694624E-4   -3.235800E-5   -3.694619E-4   -3.236380E-5   3.708767E-4   -1.749947E+2   -1.749938E+2   
7.428600E+3   2.043578E+1   2.043578E+1   -1.918000E+3   -1.918000E+3   9.000000E-4   -1.917000E+3   -1.917000E+3   -1.418286E-1   -2.038127E-1   -3.746153E-4   -3.468150E-5   -3.746148E-4   -3.468738E-5   3.762173E-4   -1.747107E+2   -1.747098E+2   
7.455548E+3   2.041189E+1   2.041189E+1   -1.928000E+3   -1.928000E+3   9.000000E-4   -1.927000E+3   -1.927000E+3   -1.395342E-1   -2.037472E-1   -3.736392E-4   -3.315627E-5   -3.736387E-4   -3.316214E-5   3.751074E-4   -1.749289E+2   -1.749280E+2   
7.483255E+3   2.041821E+1   2.041821E+1   -1.938000E+3   -1.938000E+3   9.000000E-4   -1.937000E+3   -1.937000E+3   -1.358183E-1   -2.044508E-1   -3.722165E-4   -3.020694E-5   -3.722160E-4   -3.021279E-5   3.734402E-4   -1.753604E+2   -1.753595E+2   
7.511488E+3   2.041491E+1   2.041491E+1   -1.948000E+3   -1.948000E+3   9.000000E-4   -1.947000E+3   -1.947000E+3   -1.358769E-1   -1.916886E-1   -3.639458E-4   -3.809800E-5   -3.639452E-4   -3.810372E-5   3.659345E-4   -1.740240E+2   -1.740231E+2   
7.538476E+3   2.042541E+1   2.042541E+1   -1.958000E+3   -1.958000E+3   9.000000E-4   -1.957000E+3   -1.957000E+3   -1.358064E-1   -1.972394E-1   -3.684643E-4   -3.458650E-5   -3.684637E-4   -3.459229E-5   3.700840E-4   -1.746376E+2   -1.746367E+2   
7.565426E+3   2.042510E+1   2.042510E+1   -1.968000E+3   -1.968000E+3   9.000000E-4   -1.967000E+3   -1.967000E+3   -1.421123E-1   -2.049989E-1   -3.789655E-4   -3.396596E-5   -3.789650E-4   -3.397192E-5   3.804846E-4   -1.748784E+2   -1.748775E+2   
7.593723E+3   2.041671E+1   2.041671E+1   -1.978000E+3   -1.978000E+3   9.000000E-4   -1.977000E+3   -1.977000E+3   -1.384911E-1   -2.099503E-1   -3.805958E-4   -2.845507E-5   -3.805954E-4   -2.846105E-5   3.816581E-4   -1.757243E+2   -1.757234E+2   
7.621994E+3   2.041131E+1   2.041131E+1   -1.988000E+3   -1.988000E+3   9.000000E-4   -1.988000E+3   -1.988000E+3   -1.401154E-1   -1.960690E-1   -3.726922E-4   -3.807922E-5   -3.726916E-4   -3.808507E-5   3.746325E-4   -1.741661E+2   -1.741652E+2   
7.649951E+3   2.044439E+1   2.044439E+1   -1.998000E+3   -1.998000E+3   9.000000E-4   -1.997000E+3   -1.997000E+3   -1.408019E-1   -2.103668E-1   -3.838216E-4   -2.967126E-5   -3.838211E-4   -2.967729E-5   3.849667E-4   -1.755796E+2   -1.755787E+2   
7.689981E+3   2.041760E+1   2.041760E+1   -2.098000E+3   -2.098000E+3   9.000000E-4   -2.097000E+3   -2.097000E+3   -1.410096E-1   -2.089835E-1   -3.896307E-4   -3.032100E-5   -3.896302E-4   -3.032713E-5   3.908087E-4   -1.755502E+2   -1.755493E+2   
7.718832E+3   2.043569E+1   2.043569E+1   -2.198000E+3   -2.198000E+3   9.000000E-4   -2.197000E+3   -2.197000E+3   -1.406960E-1   -2.101885E-1   -3.968981E-4   -2.902341E-5   -3.968976E-4   -2.902964E-5   3.979579E-4   -1.758177E+2   -1.758168E+2   
7.747774E+3   2.043691E+1   2.043691E+1   -2.298000E+3   -2.298000E+3   9.000000E-4   -2.298000E+3   -2.298000E+3   -1.367121E-1   -2.081053E-1   -3.993696E-4   -2.730462E-5   -3.993692E-4   -2.731090E-5   4.003020E-4   -1.760888E+2   -1.760879E+2   
7.777479E+3   2.043578E+1   2.043578E+1   -2.399000E+3   -2.399000E+3   9.000000E-4   -2.398000E+3   -2.398000E+3   -1.351201E-1   -2.045793E-1   -4.024217E-4   -2.807722E-5   -4.024213E-4   -2.808354E-5   4.034000E-4   -1.760089E+2   -1.760080E+2   
7.805921E+3   2.044052E+1   2.044052E+1   -2.499000E+3   -2.499000E+3   9.000000E-4   -2.498000E+3   -2.498000E+3   -1.309856E-1   -2.009119E-1   -4.036083E-4   -2.724033E-5   -4.036078E-4   -2.724667E-5   4.045265E-4   -1.761388E+2   -1.761379E+2   
7.834324E+3   2.043621E+1   2.043621E+1   -2.599000E+3   -2.599000E+3   9.000000E-4   -2.598000E+3   -2.598000E+3   -1.282156E-1   -1.951938E-1   -4.043004E-4   -2.858133E-5   -4.043000E-4   -2.858768E-5   4.053094E-4   -1.759563E+2   -1.759554E+2   
7.863937E+3   2.045001E+1   2.045001E+1   -2.699000E+3   -2.699000E+3   9.000000E-4   -2.698000E+3   -2.698000E+3   -1.255842E-1   -1.911811E-1   -4.062882E-4   -2.896103E-5   -4.062878E-4   -2.896741E-5   4.073191E-4   -1.759227E+2   -1.759218E+2   
7.892336E+3   2.044491E+1   2.044491E+1   -2.799000E+3   -2.799000E+3   9.000000E-4   -2.798000E+3   -2.798000E+3   -1.194049E-1   -1.889451E-1   -4.070609E-4   -2.587481E-5   -4.070605E-4   -2.588120E-5   4.078825E-4   -1.763629E+2   -1.763620E+2   
7.921208E+3   2.044698E+1   2.044698E+1   -2.899000E+3   -2.899000E+3   9.000000E-4   -2.898000E+3   -2.898000E+3   -1.181630E-1   -1.833685E-1   -4.089141E-4   -2.814826E-5   -4.089136E-4   -2.815468E-5   4.098818E-4   -1.760622E+2   -1.760613E+2   
7.950916E+3   2.043691E+1   2.043691E+1   -2.999000E+3   -2.999000E+3   9.000000E-4   -2.998000E+3   -2.998000E+3   -1.122076E-1   -1.797340E-1   -4.088588E-4   -2.607573E-5   -4.088584E-4   -2.608215E-5   4.096895E-4   -1.763508E+2   -1.763499E+2   
7.979823E+3   2.044009E+1   2.044009E+1   -3.098000E+3   -3.098000E+3   9.000000E-4   -3.098000E+3   -3.098000E+3   -1.083885E-1   -1.749657E-1   -4.094902E-4   -2.612961E-5   -4.094898E-4   -2.613605E-5   4.103230E-4   -1.763489E+2   -1.763480E+2   
8.008677E+3   2.044189E+1   2.044189E+1   -3.198000E+3   -3.198000E+3   9.000000E-4   -3.197000E+3   -3.197000E+3   -1.050468E-1   -1.695728E-1   -4.099476E-4   -2.689155E-5   -4.099472E-4   -2.689799E-5   4.108286E-4   -1.762469E+2   -1.762460E+2   
8.038424E+3   2.045760E+1   2.045760E+1   -3.298000E+3   -3.298000E+3   9.000000E-4   -3.298000E+3   -3.298000E+3   -1.001968E-1   -1.638639E-1   -4.092677E-4   -2.683518E-5   -4.092673E-4   -2.684161E-5   4.101465E-4   -1.762486E+2   -1.762477E+2   
8.067331E+3   2.045129E+1   2.045129E+1   -3.398000E+3   -3.398000E+3   9.000000E-4   -3.398000E+3   -3.398000E+3   -9.555446E-2   -1.593150E-1   -4.094815E-4   -2.620397E-5   -4.094811E-4   -2.621041E-5   4.103191E-4   -1.763385E+2   -1.763376E+2   
8.096230E+3   2.045480E+1   2.045480E+1   -3.498000E+3   -3.498000E+3   9.000000E-4   -3.498000E+3   -3.498000E+3   -9.200313E-2   -1.541970E-1   -4.100529E-4   -2.665269E-5   -4.100525E-4   -2.665913E-5   4.109182E-4   -1.762811E+2   -1.762802E+2   
8.125381E+3   2.045889E+1   2.045889E+1   -3.598000E+3   -3.598000E+3   9.000000E-4   -3.597000E+3   -3.597000E+3   -8.782171E-2   -1.501106E-1   -4.108458E-4   -2.604676E-5   -4.108454E-4   -2.605322E-5   4.116706E-4   -1.763724E+2   -1.763715E+2   
8.153633E+3   2.045690E+1   2.045690E+1   -3.698000E+3   -3.698000E+3   9.000000E-4   -3.698000E+3   -3.698000E+3   -8.402545E-2   -1.446273E-1   -4.110566E-4   -2.655431E-5   -4.110561E-4   -2.656076E-5   4.119134E-4   -1.763038E+2   -1.763029E+2   
8.183335E+3   2.045281E+1   2.045281E+1   -3.798000E+3   -3.798000E+3   9.000000E-4   -3.797000E+3   -3.797000E+3   -8.134254E-2   -1.406446E-1   -4.129633E-4   -2.688451E-5   -4.129629E-4   -2.689100E-5   4.138375E-4   -1.762752E+2   -1.762743E+2   
8.212558E+3   2.045889E+1   2.045889E+1   -3.898000E+3   -3.898000E+3   9.000000E-4   -3.897000E+3   -3.897000E+3   -7.569825E-2   -1.353312E-1   -4.119434E-4   -2.605701E-5   -4.119430E-4   -2.606348E-5   4.127667E-4   -1.763806E+2   -1.763797E+2   
8.241785E+3   2.045651E+1   2.045651E+1   -3.998000E+3   -3.998000E+3   9.000000E-4   -3.997000E+3   -3.997000E+3   -7.305468E-2   -1.312205E-1   -4.138539E-4   -2.648911E-5   -4.138535E-4   -2.649561E-5   4.147008E-4   -1.763377E+2   -1.763368E+2   
8.270957E+3   2.046319E+1   2.046319E+1   -4.098000E+3   -4.098000E+3   9.000000E-4   -4.097000E+3   -4.097000E+3   -6.907653E-2   -1.275294E-1   -4.151323E-4   -2.577121E-5   -4.151319E-4   -2.577773E-5   4.159315E-4   -1.764477E+2   -1.764468E+2   
8.299246E+3   2.046050E+1   2.046050E+1   -4.198000E+3   -4.198000E+3   9.000000E-4   -4.197000E+3   -4.197000E+3   -6.376319E-2   -1.226810E-1   -4.146694E-4   -2.487726E-5   -4.146690E-4   -2.488377E-5   4.154149E-4   -1.765668E+2   -1.765659E+2   
8.328178E+3   2.045889E+1   2.045889E+1   -4.298000E+3   -4.298000E+3   9.000000E-4   -4.298000E+3   -4.298000E+3   -5.893916E-2   -1.171791E-1   -4.141531E-4   -2.471033E-5   -4.141527E-4   -2.471683E-5   4.148896E-4   -1.765855E+2   -1.765846E+2   
8.357116E+3   2.046649E+1   2.046649E+1   -4.398000E+3   -4.398000E+3   9.000000E-4   -4.398000E+3   -4.398000E+3   -5.574040E-2   -1.110933E-1   -4.142889E-4   -2.599235E-5   -4.142885E-4   -2.599886E-5   4.151034E-4   -1.764100E+2   -1.764091E+2   
8.386816E+3   2.045931E+1   2.045931E+1   -4.499000E+3   -4.499000E+3   9.000000E-4   -4.498000E+3   -4.498000E+3   -5.203311E-2   -1.064650E-1   -4.150963E-4   -2.603440E-5   -4.150959E-4   -2.604092E-5   4.159119E-4   -1.764112E+2   -1.764103E+2   
8.415282E+3   2.046441E+1   2.046441E+1   -4.598000E+3   -4.598000E+3   9.000000E-4   -4.598000E+3   -4.598000E+3   -4.710307E-2   -1.015952E-1   -4.148846E-4   -2.540953E-5   -4.148842E-4   -2.541604E-5   4.156619E-4   -1.764953E+2   -1.764944E+2   
8.443683E+3   2.046301E+1   2.046301E+1   -4.699000E+3   -4.699000E+3   9.000000E-4   -4.698000E+3   -4.698000E+3   -4.170927E-2   -9.686221E-2   -4.144469E-4   -2.439056E-5   -4.144465E-4   -2.439707E-5   4.151640E-4   -1.766320E+2   -1.766311E+2   
8.473344E+3   2.046121E+1   2.046121E+1   -4.799000E+3   -4.799000E+3   9.000000E-4   -4.798000E+3   -4.798000E+3   -3.876373E-2   -9.372255E-2   -4.168305E-4   -2.402107E-5   -4.168301E-4   -2.402762E-5   4.175220E-4   -1.767018E+2   -1.767009E+2   
8.501327E+3   2.047231E+1   2.047231E+1   -4.899000E+3   -4.899000E+3   9.000000E-4   -4.898000E+3   -4.898000E+3   -3.392201E-2   -8.857222E-2   -4.164828E-4   -2.362851E-5   -4.164824E-4   -2.363505E-5   4.171525E-4   -1.767529E+2   -1.767520E+2   
8.529816E+3   2.048940E+1   2.048940E+1   -4.999000E+3   -4.999000E+3   9.000000E-4   -4.998000E+3   -4.998000E+3   -3.013427E-2   -8.271337E-2   -4.163690E-4   -2.437721E-5   -4.163686E-4   -2.438375E-5   4.170820E-4   -1.766493E+2   -1.766484E+2   
8.558969E+3   2.050161E+1   2.050161E+1   -5.099000E+3   -5.099000E+3   9.000000E-4   -5.098000E+3   -5.098000E+3   -2.527796E-2   -7.880162E-2   -4.168822E-4   -2.320953E-5   -4.168819E-4   -2.321607E-5   4.175278E-4   -1.768134E+2   -1.768125E+2   
8.587226E+3   2.051309E+1   2.051309E+1   -5.198000E+3   -5.198000E+3   9.000000E-4   -5.198000E+3   -5.198000E+3   -1.995271E-2   -7.501145E-2   -4.171552E-4   -2.165373E-5   -4.171548E-4   -2.166028E-5   4.177168E-4   -1.770286E+2   -1.770277E+2   
8.615527E+3   2.050280E+1   2.050280E+1   -5.299000E+3   -5.299000E+3   9.000000E-4   -5.298000E+3   -5.298000E+3   -1.775461E-2   -6.840618E-2   -4.176207E-4   -2.392465E-5   -4.176204E-4   -2.393121E-5   4.183055E-4   -1.767212E+2   -1.767203E+2   
8.645227E+3   2.051422E+1   2.051422E+1   -5.398000E+3   -5.398000E+3   9.000000E-4   -5.398000E+3   -5.398000E+3   -1.331542E-2   -6.409195E-2   -4.181407E-4   -2.328407E-5   -4.181403E-4   -2.329064E-5   4.187885E-4   -1.768128E+2   -1.768119E+2   
8.673691E+3   2.051531E+1   2.051531E+1   -5.499000E+3   -5.499000E+3   9.000000E-4   -5.498000E+3   -5.498000E+3   -9.262603E-3   -5.969239E-2   -4.188690E-4   -2.295410E-5   -4.188687E-4   -2.296068E-5   4.194975E-4   -1.768633E+2   -1.768624E+2   
8.702582E+3   2.052490E+1   2.052490E+1   -5.598000E+3   -5.598000E+3   9.000000E-4   -5.598000E+3   -5.598000E+3   -6.104370E-3   -5.490613E-2   -4.199468E-4   -2.346017E-5   -4.199465E-4   -2.346676E-5   4.206016E-4   -1.768025E+2   -1.768016E+2   
8.732289E+3   2.052920E+1   2.052920E+1   -5.699000E+3   -5.699000E+3   9.000000E-4   -5.698000E+3   -5.698000E+3   -4.402898E-4   -4.980333E-2   -4.190613E-4   -2.248935E-5   -4.190610E-4   -2.249594E-5   4.196643E-4   -1.769281E+2   -1.769272E+2   
8.761273E+3   2.053799E+1   2.053799E+1   -5.799000E+3   -5.799000E+3   9.000000E-4   -5.798000E+3   -5.798000E+3   2.420239E-3   -4.402712E-2   -4.196498E-4   -2.380584E-5   -4.196494E-4   -2.381244E-5   4.203244E-4   -1.767532E+2   -1.767523E+2   
8.790180E+3   2.054540E+1   2.054540E+1   -5.898000E+3   -5.898000E+3   9.000000E-4   -5.897000E+3   -5.897000E+3   7.126643E-3   -4.077718E-2   -4.206662E-4   -2.233269E-5   -4.206658E-4   -2.233929E-5   4.212586E-4   -1.769611E+2   -1.769602E+2   
8.819916E+3   2.054189E+1   2.054189E+1   -5.998000E+3   -5.998000E+3   9.000000E-4   -5.998000E+3   -5.998000E+3   1.199394E-2   -3.664482E-2   -4.210830E-4   -2.129056E-5   -4.210827E-4   -2.129717E-5   4.216209E-4   -1.771055E+2   -1.771046E+2   
8.858939E+3   2.053851E+1   2.053851E+1   -5.899000E+3   -5.899000E+3   9.000000E-4   -5.898000E+3   -5.898000E+3   8.537414E-3   -3.877623E-2   -4.183453E-4   -2.262413E-5   -4.183450E-4   -2.263070E-5   4.189567E-4   -1.769045E+2   -1.769036E+2   
8.886175E+3   2.053149E+1   2.053149E+1   -5.798000E+3   -5.798000E+3   9.000000E-4   -5.798000E+3   -5.798000E+3   4.272816E-3   -4.541503E-2   -4.193389E-4   -2.171173E-5   -4.193386E-4   -2.171831E-5   4.199006E-4   -1.770361E+2   -1.770352E+2   
8.913384E+3   2.054312E+1   2.054312E+1   -5.699000E+3   -5.699000E+3   9.000000E-4   -5.698000E+3   -5.698000E+3   -1.319354E-3   -4.775696E-2   -4.182329E-4   -2.434060E-5   -4.182325E-4   -2.434717E-5   4.189406E-4   -1.766692E+2   -1.766683E+2   
8.940366E+3   2.055789E+1   2.055789E+1   -5.598000E+3   -5.598000E+3   9.000000E-4   -5.598000E+3   -5.598000E+3   -3.465961E-3   -5.683551E-2   -4.194709E-4   -2.050697E-5   -4.194706E-4   -2.051356E-5   4.199718E-4   -1.772012E+2   -1.772003E+2   
8.967276E+3   2.055309E+1   2.055309E+1   -5.498000E+3   -5.498000E+3   9.000000E-4   -5.498000E+3   -5.498000E+3   -9.848228E-3   -5.900681E-2   -4.187937E-4   -2.376862E-5   -4.187933E-4   -2.377520E-5   4.194676E-4   -1.767517E+2   -1.767508E+2   
8.994248E+3   2.055270E+1   2.055270E+1   -5.399000E+3   -5.399000E+3   9.000000E-4   -5.398000E+3   -5.398000E+3   -1.417924E-2   -6.342587E-2   -4.182723E-4   -2.427221E-5   -4.182720E-4   -2.427878E-5   4.189760E-4   -1.766789E+2   -1.766780E+2   
9.021162E+3   2.054150E+1   2.054150E+1   -5.299000E+3   -5.299000E+3   9.000000E-4   -5.298000E+3   -5.298000E+3   -1.535476E-2   -7.075024E-2   -4.176021E-4   -2.087443E-5   -4.176018E-4   -2.088099E-5   4.181235E-4   -1.771384E+2   -1.771375E+2   
9.048131E+3   2.054901E+1   2.054901E+1   -5.198000E+3   -5.198000E+3   9.000000E-4   -5.198000E+3   -5.198000E+3   -2.274499E-2   -7.621501E-2   -4.199413E-4   -2.277365E-5   -4.199410E-4   -2.278025E-5   4.205584E-4   -1.768959E+2   -1.768950E+2   
9.075041E+3   2.056680E+1   2.056680E+1   -5.099000E+3   -5.099000E+3   9.000000E-4   -5.098000E+3   -5.098000E+3   -2.575968E-2   -7.804873E-2   -4.166874E-4   -2.399628E-5   -4.166870E-4   -2.400283E-5   4.173778E-4   -1.767041E+2   -1.767032E+2   
9.102226E+3   2.055569E+1   2.055569E+1   -4.999000E+3   -4.999000E+3   9.000000E-4   -4.998000E+3   -4.998000E+3   -2.982928E-2   -8.483839E-2   -4.176516E-4   -2.286051E-5   -4.176512E-4   -2.286707E-5   4.182767E-4   -1.768670E+2   -1.768661E+2   
9.129426E+3   2.055999E+1   2.055999E+1   -4.899000E+3   -4.899000E+3   9.000000E-4   -4.898000E+3   -4.898000E+3   -3.410484E-2   -9.004789E-2   -4.176476E-4   -2.283865E-5   -4.176472E-4   -2.284521E-5   4.182715E-4   -1.768700E+2   -1.768691E+2   
9.156362E+3   2.055581E+1   2.055581E+1   -4.799000E+3   -4.799000E+3   9.000000E-4   -4.798000E+3   -4.798000E+3   -3.785906E-2   -9.220362E-2   -4.151338E-4   -2.435588E-5   -4.151334E-4   -2.436240E-5   4.158477E-4   -1.766423E+2   -1.766414E+2   
9.183313E+3   2.055300E+1   2.055300E+1   -4.699000E+3   -4.699000E+3   9.000000E-4   -4.698000E+3   -4.698000E+3   -4.165077E-2   -9.944488E-2   -4.162225E-4   -2.275558E-5   -4.162222E-4   -2.276212E-5   4.168441E-4   -1.768707E+2   -1.768698E+2   
9.210591E+3   2.054531E+1   2.054531E+1   -4.599000E+3   -4.599000E+3   9.000000E-4   -4.598000E+3   -4.598000E+3   -4.623954E-2   -1.051870E-1   -4.168107E-4   -2.261363E-5   -4.168103E-4   -2.262018E-5   4.174237E-4   -1.768945E+2   -1.768936E+2   
9.237587E+3   2.055471E+1   2.055471E+1   -4.499000E+3   -4.499000E+3   9.000000E-4   -4.498000E+3   -4.498000E+3   -5.101877E-2   -1.067245E-1   -4.145742E-4   -2.519699E-5   -4.145738E-4   -2.520350E-5   4.153392E-4   -1.765220E+2   -1.765211E+2   
9.264520E+3   2.055221E+1   2.055221E+1   -4.398000E+3   -4.398000E+3   9.000000E-4   -4.398000E+3   -4.398000E+3   -5.432264E-2   -1.130855E-1   -4.147050E-4   -2.381508E-5   -4.147046E-4   -2.382159E-5   4.153882E-4   -1.767133E+2   -1.767124E+2   
9.291418E+3   2.054980E+1   2.054980E+1   -4.298000E+3   -4.298000E+3   9.000000E-4   -4.298000E+3   -4.298000E+3   -5.854274E-2   -1.158607E-1   -4.129505E-4   -2.526046E-5   -4.129501E-4   -2.526694E-5   4.137224E-4   -1.764995E+2   -1.764986E+2   
9.318634E+3   2.055270E+1   2.055270E+1   -4.198000E+3   -4.198000E+3   9.000000E-4   -4.198000E+3   -4.198000E+3   -6.347096E-2   -1.217892E-1   -4.139055E-4   -2.522989E-5   -4.139051E-4   -2.523639E-5   4.146738E-4   -1.765118E+2   -1.765109E+2   
9.345838E+3   2.055691E+1   2.055691E+1   -4.098000E+3   -4.098000E+3   9.000000E-4   -4.097000E+3   -4.097000E+3   -6.734860E-2   -1.244571E-1   -4.117714E-4   -2.651641E-5   -4.117709E-4   -2.652288E-5   4.126243E-4   -1.763155E+2   -1.763146E+2   
9.373021E+3   2.054690E+1   2.054690E+1   -3.998000E+3   -3.998000E+3   9.000000E-4   -3.997000E+3   -3.997000E+3   -7.276343E-2   -1.330423E-1   -4.149328E-4   -2.516896E-5   -4.149324E-4   -2.517548E-5   4.156954E-4   -1.765288E+2   -1.765279E+2   
9.400229E+3   2.058050E+1   2.058050E+1   -3.898000E+3   -3.898000E+3   9.000000E-4   -3.897000E+3   -3.897000E+3   -7.497464E-2   -1.369806E-1   -4.126007E-4   -2.455486E-5   -4.126003E-4   -2.456134E-5   4.133307E-4   -1.765942E+2   -1.765933E+2   
9.427420E+3   2.058419E+1   2.058419E+1   -3.798000E+3   -3.798000E+3   9.000000E-4   -3.797000E+3   -3.797000E+3   -7.717364E-2   -1.419359E-1   -4.109754E-4   -2.330411E-5   -4.109750E-4   -2.331056E-5   4.116356E-4   -1.767546E+2   -1.767537E+2   
9.454637E+3   2.059850E+1   2.059850E+1   -3.698000E+3   -3.698000E+3   9.000000E-4   -3.697000E+3   -3.697000E+3   -7.904117E-2   -1.501058E-1   -4.113806E-4   -1.984570E-5   -4.113802E-4   -1.985217E-5   4.118590E-4   -1.772381E+2   -1.772372E+2   
9.481790E+3   2.060229E+1   2.060229E+1   -3.598000E+3   -3.598000E+3   9.000000E-4   -3.598000E+3   -3.598000E+3   -7.775009E-2   -1.573616E-1   -4.090150E-4   -1.484058E-5   -4.090148E-4   -1.484701E-5   4.092842E-4   -1.779220E+2   -1.779211E+2   
9.509017E+3   2.059521E+1   2.059521E+1   -3.499000E+3   -3.499000E+3   9.000000E-4   -3.498000E+3   -3.498000E+3   -9.802749E-2   -1.490820E-1   -4.106407E-4   -3.383428E-5   -4.106402E-4   -3.384073E-5   4.120322E-4   -1.752898E+2   -1.752889E+2   
9.536217E+3   2.061630E+1   2.061630E+1   -3.398000E+3   -3.398000E+3   9.000000E-4   -3.398000E+3   -3.398000E+3   -9.963837E-2   -1.621426E-1   -4.143070E-4   -2.718238E-5   -4.143066E-4   -2.718889E-5   4.151978E-4   -1.762462E+2   -1.762453E+2   
9.563417E+3   2.060769E+1   2.060769E+1   -3.299000E+3   -3.299000E+3   9.000000E-4   -3.298000E+3   -3.298000E+3   -9.785886E-2   -1.691825E-1   -4.113839E-4   -2.198815E-5   -4.113836E-4   -2.199461E-5   4.119711E-4   -1.769405E+2   -1.769396E+2   
9.590627E+3   2.059750E+1   2.059750E+1   -3.198000E+3   -3.198000E+3   9.000000E-4   -3.198000E+3   -3.198000E+3   -1.014461E-1   -1.692906E-1   -4.073142E-4   -2.465922E-5   -4.073138E-4   -2.466562E-5   4.080600E-4   -1.765355E+2   -1.765346E+2   
9.617589E+3   2.061190E+1   2.061190E+1   -3.098000E+3   -3.098000E+3   9.000000E-4   -3.098000E+3   -3.098000E+3   -1.069564E-1   -1.741241E-1   -4.079035E-4   -2.569383E-5   -4.079031E-4   -2.570024E-5   4.087119E-4   -1.763957E+2   -1.763948E+2   
9.644729E+3   2.060491E+1   2.060491E+1   -2.999000E+3   -2.999000E+3   9.000000E-4   -2.998000E+3   -2.998000E+3   -1.106375E-1   -1.794442E-1   -4.075643E-4   -2.520685E-5   -4.075639E-4   -2.521325E-5   4.083431E-4   -1.764609E+2   -1.764600E+2   
9.671921E+3   2.060800E+1   2.060800E+1   -2.898000E+3   -2.898000E+3   9.000000E-4   -2.898000E+3   -2.898000E+3   -1.164594E-1   -1.826813E-1   -4.072474E-4   -2.743587E-5   -4.072470E-4   -2.744227E-5   4.081706E-4   -1.761459E+2   -1.761450E+2   
9.699163E+3   2.060620E+1   2.060620E+1   -2.799000E+3   -2.799000E+3   9.000000E-4   -2.798000E+3   -2.798000E+3   -1.197904E-1   -1.862619E-1   -4.054417E-4   -2.779017E-5   -4.054412E-4   -2.779654E-5   4.063930E-4   -1.760789E+2   -1.760780E+2   
9.726380E+3   2.060781E+1   2.060781E+1   -2.699000E+3   -2.699000E+3   9.000000E-4   -2.698000E+3   -2.698000E+3   -1.230101E-1   -1.925955E-1   -4.054948E-4   -2.636901E-5   -4.054943E-4   -2.637538E-5   4.063512E-4   -1.762793E+2   -1.762784E+2   
9.753559E+3   2.061910E+1   2.061910E+1   -2.599000E+3   -2.599000E+3   9.000000E-4   -2.598000E+3   -2.598000E+3   -1.246335E-1   -1.978758E-1   -4.036982E-4   -2.453326E-5   -4.036978E-4   -2.453960E-5   4.044430E-4   -1.765223E+2   -1.765214E+2   
9.780779E+3   2.061169E+1   2.061169E+1   -2.499000E+3   -2.499000E+3   9.000000E-4   -2.498000E+3   -2.498000E+3   -1.285819E-1   -2.014043E-1   -4.022847E-4   -2.533172E-5   -4.022843E-4   -2.533804E-5   4.030815E-4   -1.763969E+2   -1.763960E+2   
9.807970E+3   2.062121E+1   2.062121E+1   -2.399000E+3   -2.399000E+3   9.000000E-4   -2.398000E+3   -2.398000E+3   -1.305861E-1   -2.062817E-1   -4.004694E-4   -2.399919E-5   -4.004690E-4   -2.400548E-5   4.011878E-4   -1.765705E+2   -1.765696E+2   
9.835162E+3   2.062328E+1   2.062328E+1   -2.299000E+3   -2.299000E+3   9.000000E-4   -2.298000E+3   -2.298000E+3   -1.357740E-1   -2.063304E-1   -3.974697E-4   -2.777523E-5   -3.974693E-4   -2.778147E-5   3.984390E-4   -1.760027E+2   -1.760018E+2   
9.862377E+3   2.061929E+1   2.061929E+1   -2.198000E+3   -2.198000E+3   9.000000E-4   -2.198000E+3   -2.198000E+3   -1.373559E-1   -2.126386E-1   -3.963672E-4   -2.527667E-5   -3.963668E-4   -2.528289E-5   3.971724E-4   -1.763511E+2   -1.763502E+2   
9.889598E+3   2.062371E+1   2.062371E+1   -2.098000E+3   -2.098000E+3   9.000000E-4   -2.098000E+3   -2.098000E+3   -1.381055E-1   -2.121255E-1   -3.898894E-4   -2.643770E-5   -3.898889E-4   -2.644382E-5   3.907847E-4   -1.761208E+2   -1.761199E+2   
9.916757E+3   2.062280E+1   2.062280E+1   -1.998000E+3   -1.998000E+3   9.000000E-4   -1.998000E+3   -1.998000E+3   -1.391455E-1   -2.052768E-1   -3.791576E-4   -3.170755E-5   -3.791571E-4   -3.171351E-5   3.804811E-4   -1.752197E+2   -1.752188E+2   
9.955544E+3   2.061740E+1   2.061740E+1   -1.948000E+3   -1.948000E+3   9.000000E-4   -1.948000E+3   -1.948000E+3   -1.364105E-1   -2.048679E-1   -3.736513E-4   -3.030666E-5   -3.736508E-4   -3.031253E-5   3.748784E-4   -1.753629E+2   -1.753620E+2   
9.982495E+3   2.060940E+1   2.060940E+1   -1.898000E+3   -1.898000E+3   9.000000E-4   -1.898000E+3   -1.898000E+3   -1.355171E-1   -2.051275E-1   -3.698944E-4   -2.972179E-5   -3.698939E-4   -2.972760E-5   3.710866E-4   -1.754060E+2   -1.754051E+2   
1.000949E+4   2.059969E+1   2.059969E+1   -1.849000E+3   -1.849000E+3   9.000000E-4   -1.847000E+3   -1.847000E+3   -1.341508E-1   -2.026432E-1   -3.638129E-4   -3.052033E-5   -3.638125E-4   -3.052604E-5   3.650909E-4   -1.752047E+2   -1.752038E+2   
1.003639E+4   2.061599E+1   2.061599E+1   -1.798000E+3   -1.798000E+3   9.000000E-4   -1.798000E+3   -1.798000E+3   -1.334857E-1   -2.009540E-1   -3.589104E-4   -3.128864E-5   -3.589099E-4   -3.129428E-5   3.602717E-4   -1.750177E+2   -1.750168E+2   
1.006330E+4   2.061770E+1   2.061770E+1   -1.748000E+3   -1.748000E+3   9.000000E-4   -1.748000E+3   -1.748000E+3   -1.338117E-1   -1.967118E-1   -3.528347E-4   -3.429944E-5   -3.528342E-4   -3.430498E-5   3.544980E-4   -1.744477E+2   -1.744468E+2   
1.009026E+4   2.062731E+1   2.062731E+1   -1.698000E+3   -1.698000E+3   9.000000E-4   -1.698000E+3   -1.698000E+3   -1.327446E-1   -1.978959E-1   -3.496073E-4   -3.302739E-5   -3.496068E-4   -3.303288E-5   3.511639E-4   -1.746033E+2   -1.746024E+2   
1.011719E+4   2.064019E+1   2.064019E+1   -1.649000E+3   -1.649000E+3   9.000000E-4   -1.648000E+3   -1.648000E+3   -1.299837E-1   -1.975113E-1   -3.441001E-4   -3.159417E-5   -3.440996E-4   -3.159958E-5   3.455475E-4   -1.747540E+2   -1.747531E+2   
1.014413E+4   2.064321E+1   2.064321E+1   -1.598000E+3   -1.598000E+3   9.000000E-4   -1.597000E+3   -1.597000E+3   -1.290361E-1   -1.920285E-1   -3.362007E-4   -3.452506E-5   -3.362002E-4   -3.453034E-5   3.379688E-4   -1.741367E+2   -1.741358E+2   
1.017108E+4   2.065469E+1   2.065469E+1   -1.548000E+3   -1.548000E+3   9.000000E-4   -1.548000E+3   -1.548000E+3   -1.274173E-1   -1.912023E-1   -3.312427E-4   -3.412349E-5   -3.312421E-4   -3.412869E-5   3.329957E-4   -1.741183E+2   -1.741174E+2   
1.019798E+4   2.066061E+1   2.066061E+1   -1.499000E+3   -1.499000E+3   9.000000E-4   -1.498000E+3   -1.498000E+3   -1.280486E-1   -1.859959E-1   -3.247009E-4   -3.793398E-5   -3.247003E-4   -3.793908E-5   3.269092E-4   -1.733365E+2   -1.733356E+2   
1.022516E+4   2.064910E+1   2.064910E+1   -1.449000E+3   -1.449000E+3   9.000000E-4   -1.448000E+3   -1.448000E+3   -1.250930E-1   -1.875060E-1   -3.203909E-4   -3.519998E-5   -3.203904E-4   -3.520501E-5   3.223187E-4   -1.737303E+2   -1.737294E+2   
1.025215E+4   2.066271E+1   2.066271E+1   -1.399000E+3   -1.399000E+3   9.000000E-4   -1.398000E+3   -1.398000E+3   -1.233389E-1   -1.843054E-1   -3.136026E-4   -3.617882E-5   -3.136021E-4   -3.618375E-5   3.156826E-4   -1.734192E+2   -1.734183E+2   
1.027908E+4   2.065859E+1   2.065859E+1   -1.349000E+3   -1.349000E+3   9.000000E-4   -1.349000E+3   -1.349000E+3   -1.222234E-1   -1.829297E-1   -3.086077E-4   -3.645282E-5   -3.086072E-4   -3.645767E-5   3.107532E-4   -1.732634E+2   -1.732625E+2   
1.030623E+4   2.065939E+1   2.065939E+1   -1.299000E+3   -1.299000E+3   9.000000E-4   -1.299000E+3   -1.299000E+3   -1.203927E-1   -1.810936E-1   -3.027259E-4   -3.653746E-5   -3.027253E-4   -3.654221E-5   3.049229E-4   -1.731180E+2   -1.731171E+2   
1.033344E+4   2.065701E+1   2.065701E+1   -1.249000E+3   -1.249000E+3   9.000000E-4   -1.248000E+3   -1.248000E+3   -1.182577E-1   -1.771559E-1   -2.950883E-4   -3.772099E-5   -2.950877E-4   -3.772563E-5   2.974895E-4   -1.727154E+2   -1.727145E+2   
1.036042E+4   2.065331E+1   2.065331E+1   -1.199000E+3   -1.199000E+3   9.000000E-4   -1.199000E+3   -1.199000E+3   -1.171054E-1   -1.732874E-1   -2.883148E-4   -3.951076E-5   -2.883142E-4   -3.951529E-5   2.910095E-4   -1.721968E+2   -1.721959E+2   
1.038760E+4   2.066000E+1   2.066000E+1   -1.149000E+3   -1.149000E+3   9.000000E-4   -1.148000E+3   -1.148000E+3   -1.140687E-1   -1.705171E-1   -2.808718E-4   -3.937121E-5   -2.808712E-4   -3.937562E-5   2.836178E-4   -1.720206E+2   -1.720197E+2   
1.041478E+4   2.065359E+1   2.065359E+1   -1.099000E+3   -1.099000E+3   9.000000E-4   -1.099000E+3   -1.099000E+3   -1.117631E-1   -1.689957E-1   -2.749477E-4   -3.894086E-5   -2.749471E-4   -3.894518E-5   2.776916E-4   -1.719388E+2   -1.719379E+2   
1.044174E+4   2.064239E+1   2.064239E+1   -1.049000E+3   -1.049000E+3   9.000000E-4   -1.049000E+3   -1.049000E+3   -1.111723E-1   -1.646086E-1   -2.681332E-4   -4.142934E-5   -2.681325E-4   -4.143355E-5   2.713149E-4   -1.712167E+2   -1.712158E+2   
1.046889E+4   2.064791E+1   2.064791E+1   -1.000000E+3   -1.000000E+3   9.000000E-4   -9.990000E+2   -9.990000E+2   -1.064135E-1   -1.644071E-1   -2.613669E-4   -3.854951E-5   -2.613663E-4   -3.855362E-5   2.641945E-4   -1.716098E+2   -1.716089E+2   
1.049569E+4   2.063870E+1   2.063870E+1   -9.490000E+2   -9.490000E+2   9.000000E-4   -9.490000E+2   -9.490000E+2   -1.053800E-1   -1.595850E-1   -2.539388E-4   -4.101134E-5   -2.539382E-4   -4.101533E-5   2.572292E-4   -1.708259E+2   -1.708250E+2   
1.052249E+4   2.065261E+1   2.065261E+1   -8.990000E+2   -8.990000E+2   9.000000E-4   -8.990000E+2   -8.990000E+2   -1.019061E-1   -1.556559E-1   -2.454436E-4   -4.129254E-5   -2.454429E-4   -4.129640E-5   2.488928E-4   -1.704502E+2   -1.704493E+2   
1.054933E+4   2.065051E+1   2.065051E+1   -8.490000E+2   -8.490000E+2   9.000000E-4   -8.490000E+2   -8.490000E+2   -9.809266E-2   -1.524175E-1   -2.371983E-4   -4.092029E-5   -2.371976E-4   -4.092402E-5   2.407021E-4   -1.702120E+2   -1.702111E+2   
1.057611E+4   2.064440E+1   2.064440E+1   -7.990000E+2   -7.990000E+2   9.000000E-4   -7.990000E+2   -7.990000E+2   -9.605569E-2   -1.476045E-1   -2.290796E-4   -4.270676E-5   -2.290789E-4   -4.271035E-5   2.330265E-4   -1.694397E+2   -1.694388E+2   
1.060292E+4   2.063400E+1   2.063400E+1   -7.500000E+2   -7.500000E+2   9.000000E-4   -7.490000E+2   -7.490000E+2   -9.192970E-2   -1.453781E-1   -2.213288E-4   -4.150059E-5   -2.213281E-4   -4.150407E-5   2.251860E-4   -1.693800E+2   -1.693791E+2   
1.062970E+4   2.065151E+1   2.065151E+1   -6.990000E+2   -6.990000E+2   9.000000E-4   -6.990000E+2   -6.990000E+2   -8.884092E-2   -1.396576E-1   -2.118413E-4   -4.314575E-5   -2.118406E-4   -4.314908E-5   2.161904E-4   -1.684880E+2   -1.684871E+2   
1.065656E+4   2.064919E+1   2.064919E+1   -6.490000E+2   -6.490000E+2   9.000000E-4   -6.490000E+2   -6.490000E+2   -8.467865E-2   -1.360229E-1   -2.030749E-4   -4.278563E-5   -2.030742E-4   -4.278882E-5   2.075332E-4   -1.681024E+2   -1.681015E+2   
1.068332E+4   2.063979E+1   2.063979E+1   -5.990000E+2   -5.990000E+2   9.000000E-4   -5.990000E+2   -5.990000E+2   -7.969560E-2   -1.297565E-1   -1.918875E-4   -4.350390E-5   -1.918868E-4   -4.350691E-5   1.967572E-4   -1.672261E+2   -1.672252E+2   
1.071010E+4   2.063439E+1   2.063439E+1   -5.490000E+2   -5.490000E+2   9.000000E-4   -5.490000E+2   -5.490000E+2   -8.173890E-2   -1.217596E-1   -1.843642E-4   -4.998106E-5   -1.843634E-4   -4.998396E-5   1.910190E-4   -1.648317E+2   -1.648308E+2   
1.073689E+4   2.062951E+1   2.062951E+1   -4.990000E+2   -4.990000E+2   9.000000E-4   -4.980000E+2   -4.980000E+2   -6.782422E-2   -1.241698E-1   -1.730078E-4   -3.937992E-5   -1.730072E-4   -3.938264E-5   1.774331E-4   -1.671769E+2   -1.671760E+2   
1.076373E+4   2.062261E+1   2.062261E+1   -4.490000E+2   -4.490000E+2   9.000000E-4   -4.480000E+2   -4.480000E+2   -6.522359E-2   -1.148046E-1   -1.612962E-4   -4.360317E-5   -1.612956E-4   -4.360570E-5   1.670859E-4   -1.648728E+2   -1.648719E+2   
1.079052E+4   2.062991E+1   2.062991E+1   -3.990000E+2   -3.990000E+2   9.000000E-4   -3.980000E+2   -3.980000E+2   -5.934566E-2   -1.121509E-1   -1.520280E-4   -4.149168E-5   -1.520273E-4   -4.149406E-5   1.575883E-4   -1.647345E+2   -1.647336E+2   
1.081732E+4   2.063580E+1   2.063580E+1   -3.490000E+2   -3.490000E+2   9.000000E-4   -3.480000E+2   -3.480000E+2   -5.172999E-2   -1.045499E-1   -1.380732E-4   -4.127758E-5   -1.380726E-4   -4.127975E-5   1.441113E-4   -1.633557E+2   -1.633548E+2   
1.084410E+4   2.063940E+1   2.063940E+1   -2.990000E+2   -2.990000E+2   9.000000E-4   -2.980000E+2   -2.980000E+2   -4.373152E-2   -9.495660E-2   -1.224515E-4   -4.203908E-5   -1.224509E-4   -4.204100E-5   1.294668E-4   -1.610520E+2   -1.610511E+2   
1.087091E+4   2.064919E+1   2.064919E+1   -2.490000E+2   -2.490000E+2   9.000000E-4   -2.480000E+2   -2.480000E+2   -3.625844E-2   -9.345322E-2   -1.128841E-4   -3.815215E-5   -1.128835E-4   -3.815392E-5   1.191570E-4   -1.613260E+2   -1.613251E+2   
1.089772E+4   2.065151E+1   2.065151E+1   -1.990000E+2   -1.990000E+2   9.000000E-4   -1.980000E+2   -1.980000E+2   -3.026653E-2   -7.445995E-2   -9.204562E-5   -4.606152E-5   -9.204490E-5   -4.606297E-5   1.029275E-4   -1.534157E+2   -1.534148E+2   
1.092452E+4   2.064761E+1   2.064761E+1   -1.490000E+2   -1.490000E+2   9.000000E-4   -1.480000E+2   -1.480000E+2   -2.088630E-2   -6.576261E-2   -7.609412E-5   -4.534714E-5   -7.609341E-5   -4.534834E-5   8.858148E-5   -1.492078E+2   -1.492069E+2   
1.095127E+4   2.063979E+1   2.063979E+1   -9.900000E+1   -9.900000E+1   9.000000E-4   -9.800000E+1   -9.800000E+1   -6.671419E-3   -6.738452E-2   -6.404125E-5   -3.502930E-5   -6.404070E-5   -3.503030E-5   7.299543E-5   -1.513222E+2   -1.513213E+2   
1.097786E+4   2.063500E+1   2.063500E+1   -4.900000E+1   -4.900000E+1   9.000000E-4   -4.900000E+1   -4.900000E+1   7.283255E-3   -4.490222E-2   -3.528401E-5   -3.977666E-5   -3.528338E-5   -3.977721E-5   5.317089E-5   -1.315747E+2   -1.315738E+2   
1.100438E+4   2.065511E+1   2.065511E+1   0.000000E+0   0.000000E+0   9.000000E-4   0.000000E+0   0.000000E+0   2.812177E-2   -2.487484E-2   -3.471224E-6   -3.841254E-5   -3.470621E-6   -3.841259E-5   3.856906E-5   -9.516362E+1   -9.516272E+1   
1.104270E+4   2.065139E+1   2.065139E+1   9.000000E+0   9.000000E+0   9.000000E-4   1.000000E+1   1.000000E+1   3.046732E-2   -1.686853E-2   4.452444E-6   -4.182883E-5   4.453101E-6   -4.182876E-5   4.206513E-5   -8.392407E+1   -8.392317E+1   
1.106949E+4   2.064999E+1   2.064999E+1   1.900000E+1   1.900000E+1   9.000000E-4   2.000000E+1   2.000000E+1   3.643364E-2   -1.922630E-2   7.602709E-6   -3.642413E-5   7.603281E-6   -3.642401E-5   3.720912E-5   -7.821008E+1   -7.820918E+1   
1.109632E+4   2.063741E+1   2.063741E+1   2.900000E+1   2.900000E+1   9.000000E-4   3.000000E+1   3.000000E+1   3.942640E-2   -1.507964E-2   1.326163E-5   -3.702344E-5   1.326222E-5   -3.702323E-5   3.932691E-5   -7.029270E+1   -7.029180E+1   
1.112313E+4   2.065090E+1   2.065090E+1   3.900000E+1   3.900000E+1   9.000000E-4   4.000000E+1   4.000000E+1   4.258736E-2   -6.813413E-3   2.193452E-5   -4.005612E-5   2.193515E-5   -4.005578E-5   4.566855E-5   -6.129512E+1   -6.129422E+1   
1.114992E+4   2.064459E+1   2.064459E+1   4.900000E+1   4.900000E+1   9.000000E-4   5.000000E+1   5.000000E+1   4.724931E-2   -6.720784E-3   2.590195E-5   -3.703620E-5   2.590254E-5   -3.703579E-5   4.519504E-5   -5.503227E+1   -5.503137E+1   
1.117668E+4   2.064019E+1   2.064019E+1   5.900000E+1   5.900000E+1   9.000000E-4   6.000000E+1   6.000000E+1   5.011294E-2   -3.060413E-3   3.112918E-5   -3.742119E-5   3.112977E-5   -3.742070E-5   4.867619E-5   -5.024429E+1   -5.024339E+1   
1.120353E+4   2.065960E+1   2.065960E+1   6.900000E+1   6.900000E+1   9.000000E-4   7.000000E+1   7.000000E+1   5.251887E-2   1.322706E-3   3.654675E-5   -3.855827E-5   3.654736E-5   -3.855770E-5   5.312632E-5   -4.653417E+1   -4.653327E+1   
1.123032E+4   2.065670E+1   2.065670E+1   7.900000E+1   7.900000E+1   9.000000E-4   8.000000E+1   8.000000E+1   5.636449E-2   4.239303E-3   4.193308E-5   -3.782824E-5   4.193367E-5   -3.782758E-5   5.647441E-5   -4.205393E+1   -4.205303E+1   
1.125712E+4   2.065759E+1   2.065759E+1   8.900000E+1   8.900000E+1   9.000000E-4   9.000000E+1   9.000000E+1   5.981732E-2   2.560097E-3   4.381451E-5   -3.452044E-5   4.381505E-5   -3.451975E-5   5.577967E-5   -3.823376E+1   -3.823286E+1   
1.128394E+4   2.063690E+1   2.063690E+1   9.900000E+1   9.900000E+1   9.000000E-4   1.000000E+2   1.000000E+2   6.025731E-2   1.087263E-2   5.062979E-5   -3.939779E-5   5.063041E-5   -3.939700E-5   6.415265E-5   -3.788842E+1   -3.788752E+1   
1.131096E+4   2.064611E+1   2.064611E+1   1.090000E+2   1.090000E+2   9.000000E-4   1.100000E+2   1.100000E+2   6.448591E-2   1.206127E-2   5.506696E-5   -3.734438E-5   5.506755E-5   -3.734351E-5   6.653550E-5   -3.414367E+1   -3.414277E+1   
1.133797E+4   2.064321E+1   2.064321E+1   1.190000E+2   1.190000E+2   9.000000E-4   1.200000E+2   1.200000E+2   6.772884E-2   1.155151E-2   5.762500E-5   -3.489931E-5   5.762555E-5   -3.489841E-5   6.736915E-5   -3.120027E+1   -3.119937E+1   
1.136501E+4   2.065069E+1   2.065069E+1   1.290000E+2   1.290000E+2   9.000000E-4   1.300000E+2   1.300000E+2   6.932637E-2   1.567777E-2   6.230036E-5   -3.641722E-5   6.230093E-5   -3.641624E-5   7.216335E-5   -3.030811E+1   -3.030721E+1   
1.139200E+4   2.064889E+1   2.064889E+1   1.390000E+2   1.390000E+2   9.000000E-4   1.400000E+2   1.400000E+2   7.172983E-2   1.678352E-2   6.541137E-5   -3.553073E-5   6.541193E-5   -3.552971E-5   7.443844E-5   -2.851032E+1   -2.850942E+1   
1.141902E+4   2.064831E+1   2.064831E+1   1.490000E+2   1.490000E+2   9.000000E-4   1.490000E+2   1.490000E+2   7.246292E-2   1.925983E-2   6.825951E-5   -3.660259E-5   6.826008E-5   -3.660152E-5   7.745392E-5   -2.820141E+1   -2.820051E+1   
1.144597E+4   2.064739E+1   2.064739E+1   1.590000E+2   1.590000E+2   9.000000E-4   1.600000E+2   1.600000E+2   7.552089E-2   1.878662E-2   7.078115E-5   -3.430700E-5   7.078169E-5   -3.430588E-5   7.865711E-5   -2.585906E+1   -2.585816E+1   
1.147307E+4   2.064059E+1   2.064059E+1   1.690000E+2   1.690000E+2   9.000000E-4   1.700000E+2   1.700000E+2   7.727871E-2   2.381903E-2   7.620511E-5   -3.627787E-5   7.620568E-5   -3.627668E-5   8.439966E-5   -2.545705E+1   -2.545615E+1   
1.150008E+4   2.063931E+1   2.063931E+1   1.790000E+2   1.790000E+2   9.000000E-4   1.800000E+2   1.800000E+2   7.906943E-2   2.390284E-2   7.817178E-5   -3.516885E-5   7.817233E-5   -3.516763E-5   8.571858E-5   -2.422260E+1   -2.422170E+1   
1.152717E+4   2.064581E+1   2.064581E+1   1.890000E+2   1.890000E+2   9.000000E-4   1.900000E+2   1.900000E+2   8.117490E-2   2.754676E-2   8.286077E-5   -3.604969E-5   8.286134E-5   -3.604839E-5   9.036309E-5   -2.351210E+1   -2.351120E+1   
1.155418E+4   2.064480E+1   2.064480E+1   1.990000E+2   1.990000E+2   9.000000E-4   2.000000E+2   2.000000E+2   8.218071E-2   2.485960E-2   8.233348E-5   -3.375225E-5   8.233401E-5   -3.375095E-5   8.898323E-5   -2.229096E+1   -2.229006E+1   
1.158108E+4   2.064001E+1   2.064001E+1   2.090000E+2   2.090000E+2   9.000000E-4   2.100000E+2   2.100000E+2   8.448516E-2   2.958398E-2   8.792054E-5   -3.516794E-5   8.792110E-5   -3.516655E-5   9.469322E-5   -2.180125E+1   -2.180035E+1   
1.160810E+4   2.063629E+1   2.063629E+1   2.190000E+2   2.190000E+2   9.000000E-4   2.200000E+2   2.200000E+2   8.568357E-2   3.030003E-2   8.992039E-5   -3.484492E-5   8.992094E-5   -3.484351E-5   9.643570E-5   -2.118178E+1   -2.118088E+1   
1.163514E+4   2.064440E+1   2.064440E+1   2.290000E+2   2.290000E+2   9.000000E-4   2.300000E+2   2.300000E+2   8.803921E-2   3.383306E-2   9.470518E-5   -3.549026E-5   9.470574E-5   -3.548878E-5   1.011367E-4   -2.054322E+1   -2.054232E+1   
1.166212E+4   2.062679E+1   2.062679E+1   2.390000E+2   2.390000E+2   9.000000E-4   2.400000E+2   2.400000E+2   8.918217E-2   3.472552E-2   9.679057E-5   -3.531328E-5   9.679112E-5   -3.531176E-5   1.030313E-4   -2.004410E+1   -2.004320E+1   
1.168912E+4   2.062499E+1   2.062499E+1   2.490000E+2   2.490000E+2   9.000000E-4   2.500000E+2   2.500000E+2   8.978149E-2   3.723289E-2   9.963400E-5   -3.649705E-5   9.963457E-5   -3.649549E-5   1.061083E-4   -2.011835E+1   -2.011745E+1   
1.171613E+4   2.063561E+1   2.063561E+1   2.590000E+2   2.590000E+2   9.000000E-4   2.600000E+2   2.600000E+2   9.138791E-2   3.680846E-2   1.011152E-4   -3.519697E-5   1.011158E-4   -3.519538E-5   1.070659E-4   -1.919238E+1   -1.919148E+1   
1.174315E+4   2.063979E+1   2.063979E+1   2.690000E+2   2.690000E+2   9.000000E-4   2.700000E+2   2.700000E+2   9.466841E-2   4.053738E-2   1.066802E-4   -3.534608E-5   1.066808E-4   -3.534440E-5   1.123834E-4   -1.833144E+1   -1.833054E+1   
1.177016E+4   2.063711E+1   2.063711E+1   2.790000E+2   2.790000E+2   9.000000E-4   2.800000E+2   2.800000E+2   9.538321E-2   4.155479E-2   1.085561E-4   -3.553207E-5   1.085566E-4   -3.553036E-5   1.142232E-4   -1.812407E+1   -1.812317E+1   
1.179718E+4   2.063580E+1   2.063580E+1   2.890000E+2   2.890000E+2   9.000000E-4   2.900000E+2   2.900000E+2   9.576471E-2   4.436655E-2   1.114623E-4   -3.704931E-5   1.114628E-4   -3.704756E-5   1.174584E-4   -1.838646E+1   -1.838556E+1   
1.182421E+4   2.064510E+1   2.064510E+1   2.990000E+2   2.990000E+2   9.000000E-4   3.000000E+2   3.000000E+2   9.870572E-2   4.391468E-2   1.138513E-4   -3.484153E-5   1.138518E-4   -3.483974E-5   1.190632E-4   -1.701551E+1   -1.701461E+1   
1.185117E+4   2.065029E+1   2.065029E+1   3.090000E+2   3.090000E+2   9.000000E-4   3.100000E+2   3.100000E+2   9.916859E-2   4.713902E-2   1.171041E-4   -3.655941E-5   1.171047E-4   -3.655757E-5   1.226783E-4   -1.733814E+1   -1.733724E+1   
1.187826E+4   2.063961E+1   2.063961E+1   3.190000E+2   3.190000E+2   9.000000E-4   3.200000E+2   3.200000E+2   1.011196E-1   4.616214E-2   1.184362E-4   -3.468796E-5   1.184368E-4   -3.468610E-5   1.234115E-4   -1.632441E+1   -1.632351E+1   
1.190531E+4   2.065151E+1   2.065151E+1   3.290000E+2   3.290000E+2   9.000000E-4   3.300000E+2   3.300000E+2   1.016294E-1   4.880024E-2   1.213094E-4   -3.601229E-5   1.213099E-4   -3.601038E-5   1.265419E-4   -1.653422E+1   -1.653332E+1   
1.193234E+4   2.065359E+1   2.065359E+1   3.390000E+2   3.390000E+2   9.000000E-4   3.400000E+2   3.400000E+2   1.035417E-1   4.774628E-2   1.225603E-4   -3.411904E-5   1.225609E-4   -3.411712E-5   1.272209E-4   -1.555644E+1   -1.555554E+1   
1.195932E+4   2.065200E+1   2.065200E+1   3.490000E+2   3.490000E+2   9.000000E-4   3.500000E+2   3.500000E+2   1.037233E-1   5.095021E-2   1.256035E-4   -3.601205E-5   1.256040E-4   -3.601007E-5   1.306641E-4   -1.599824E+1   -1.599734E+1   
1.198640E+4   2.064880E+1   2.064880E+1   3.590000E+2   3.590000E+2   9.000000E-4   3.600000E+2   3.600000E+2   1.040167E-1   5.293442E-2   1.278665E-4   -3.707669E-5   1.278671E-4   -3.707468E-5   1.331335E-4   -1.617026E+1   -1.616936E+1   
1.201344E+4   2.064489E+1   2.064489E+1   3.690000E+2   3.690000E+2   9.000000E-4   3.700000E+2   3.700000E+2   1.050045E-1   5.405906E-2   1.300074E-4   -3.714671E-5   1.300080E-4   -3.714467E-5   1.352102E-4   -1.594610E+1   -1.594520E+1   
1.204049E+4   2.065060E+1   2.065060E+1   3.790000E+2   3.790000E+2   9.000000E-4   3.800000E+2   3.800000E+2   1.090244E-1   5.190818E-2   1.319511E-4   -3.316895E-5   1.319516E-4   -3.316687E-5   1.360561E-4   -1.411026E+1   -1.410936E+1   
1.206757E+4   2.065161E+1   2.065161E+1   3.890000E+2   3.890000E+2   9.000000E-4   3.890000E+2   3.890000E+2   1.098669E-1   5.636625E-2   1.362689E-4   -3.539240E-5   1.362694E-4   -3.539026E-5   1.407900E-4   -1.455944E+1   -1.455854E+1   
1.209465E+4   2.064651E+1   2.064651E+1   3.990000E+2   3.990000E+2   9.000000E-4   4.000000E+2   4.000000E+2   1.103151E-1   5.455667E-2   1.360378E-4   -3.401284E-5   1.360383E-4   -3.401071E-5   1.402253E-4   -1.403759E+1   -1.403669E+1   
1.212167E+4   2.064529E+1   2.064529E+1   4.090000E+2   4.090000E+2   9.000000E-4   4.100000E+2   4.100000E+2   1.115160E-1   5.803328E-2   1.399807E-4   -3.539408E-5   1.399812E-4   -3.539188E-5   1.443861E-4   -1.418981E+1   -1.418891E+1   
1.214863E+4   2.063171E+1   2.063171E+1   4.190000E+2   4.190000E+2   9.000000E-4   4.200000E+2   4.200000E+2   1.119626E-1   5.905158E-2   1.416709E-4   -3.575957E-5   1.416714E-4   -3.575735E-5   1.461143E-4   -1.416629E+1   -1.416539E+1   
1.217573E+4   2.065069E+1   2.065069E+1   4.290000E+2   4.290000E+2   9.000000E-4   4.290000E+2   4.290000E+2   1.126759E-1   6.170158E-2   1.446274E-4   -3.695196E-5   1.446280E-4   -3.694969E-5   1.492734E-4   -1.433232E+1   -1.433142E+1   
1.220278E+4   2.063229E+1   2.063229E+1   4.390000E+2   4.390000E+2   9.000000E-4   4.400000E+2   4.400000E+2   1.133399E-1   6.236917E-2   1.462883E-4   -3.695916E-5   1.462889E-4   -3.695687E-5   1.508849E-4   -1.417885E+1   -1.417795E+1   
1.222983E+4   2.065029E+1   2.065029E+1   4.490000E+2   4.490000E+2   9.000000E-4   4.500000E+2   4.500000E+2   1.146739E-1   6.387743E-2   1.489394E-4   -3.703520E-5   1.489400E-4   -3.703286E-5   1.534749E-4   -1.396393E+1   -1.396303E+1   
1.225690E+4   2.062100E+1   2.062100E+1   4.590000E+2   4.590000E+2   9.000000E-4   4.600000E+2   4.600000E+2   1.158082E-1   6.375435E-2   1.503047E-4   -3.623640E-5   1.503052E-4   -3.623403E-5   1.546110E-4   -1.355457E+1   -1.355367E+1   
1.228399E+4   2.062991E+1   2.062991E+1   4.690000E+2   4.690000E+2   9.000000E-4   4.690000E+2   4.690000E+2   1.171023E-1   6.380187E-2   1.518344E-4   -3.543299E-5   1.518350E-4   -3.543060E-5   1.559140E-4   -1.313580E+1   -1.313490E+1   
1.231103E+4   2.064529E+1   2.064529E+1   4.790000E+2   4.790000E+2   9.000000E-4   4.800000E+2   4.800000E+2   1.196109E-1   6.461025E-2   1.548757E-4   -3.429601E-5   1.548762E-4   -3.429358E-5   1.586276E-4   -1.248621E+1   -1.248531E+1   
1.233813E+4   2.064971E+1   2.064971E+1   4.890000E+2   4.890000E+2   9.000000E-4   4.890000E+2   4.890000E+2   1.195698E-1   6.762739E-2   1.575664E-4   -3.621881E-5   1.575669E-4   -3.621634E-5   1.616755E-4   -1.294536E+1   -1.294446E+1   
1.236518E+4   2.064160E+1   2.064160E+1   4.990000E+2   4.990000E+2   9.000000E-4   5.000000E+2   5.000000E+2   1.205530E-1   6.773005E-2   1.590517E-4   -3.566380E-5   1.590523E-4   -3.566130E-5   1.630011E-4   -1.263826E+1   -1.263736E+1   
1.239224E+4   2.064431E+1   2.064431E+1   5.090000E+2   5.090000E+2   9.000000E-4   5.100000E+2   5.100000E+2   1.202934E-1   7.053847E-2   1.615102E-4   -3.760688E-5   1.615108E-4   -3.760434E-5   1.658307E-4   -1.310749E+1   -1.310659E+1   
1.241934E+4   2.065429E+1   2.065429E+1   5.190000E+2   5.190000E+2   9.000000E-4   5.200000E+2   5.200000E+2   1.232231E-1   7.021486E-2   1.639816E-4   -3.548590E-5   1.639821E-4   -3.548333E-5   1.677773E-4   -1.221062E+1   -1.220972E+1   
1.244640E+4   2.063271E+1   2.063271E+1   5.290000E+2   5.290000E+2   9.000000E-4   5.300000E+2   5.300000E+2   1.240366E-1   7.180085E-2   1.663258E-4   -3.595734E-5   1.663264E-4   -3.595473E-5   1.701682E-4   -1.219882E+1   -1.219792E+1   
1.247344E+4   2.066589E+1   2.066589E+1   5.390000E+2   5.390000E+2   9.000000E-4   5.400000E+2   5.400000E+2   1.238030E-1   7.185841E-2   1.668678E-4   -3.618324E-5   1.668683E-4   -3.618062E-5   1.707457E-4   -1.223449E+1   -1.223359E+1   
1.250052E+4   2.065151E+1   2.065151E+1   5.480000E+2   5.480000E+2   9.000000E-4   5.490000E+2   5.490000E+2   1.244410E-1   7.523723E-2   1.702846E-4   -3.787626E-5   1.702851E-4   -3.787358E-5   1.744461E-4   -1.254011E+1   -1.253921E+1   
1.252758E+4   2.065240E+1   2.065240E+1   5.590000E+2   5.590000E+2   9.000000E-4   5.590000E+2   5.590000E+2   1.264002E-1   7.316345E-2   1.708509E-4   -3.532150E-5   1.708515E-4   -3.531882E-5   1.744639E-4   -1.168070E+1   -1.167980E+1   
1.255512E+4   2.065051E+1   2.065051E+1   5.680000E+2   5.680000E+2   9.000000E-4   5.690000E+2   5.690000E+2   1.269352E-1   7.386488E-2   1.723797E-4   -3.543220E-5   1.723802E-4   -3.542949E-5   1.759835E-4   -1.161522E+1   -1.161432E+1   
1.258260E+4   2.065811E+1   2.065811E+1   5.780000E+2   5.780000E+2   9.000000E-4   5.790000E+2   5.790000E+2   1.286013E-1   7.326582E-2   1.737795E-4   -3.398439E-5   1.737801E-4   -3.398166E-5   1.770714E-4   -1.106514E+1   -1.106424E+1   
1.261010E+4   2.067660E+1   2.067660E+1   5.880000E+2   5.880000E+2   9.000000E-4   5.890000E+2   5.890000E+2   1.280002E-1   7.717547E-2   1.767752E-4   -3.683593E-5   1.767758E-4   -3.683315E-5   1.805723E-4   -1.177070E+1   -1.176980E+1   
1.263764E+4   2.066750E+1   2.066750E+1   5.980000E+2   5.980000E+2   9.000000E-4   5.990000E+2   5.990000E+2   1.296712E-1   7.452425E-2   1.767353E-4   -3.411673E-5   1.767358E-4   -3.411395E-5   1.799981E-4   -1.092591E+1   -1.092501E+1   
1.266510E+4   2.067309E+1   2.067309E+1   6.080000E+2   6.080000E+2   9.000000E-4   6.090000E+2   6.090000E+2   1.324777E-1   7.084286E-2   1.767597E-4   -3.000303E-5   1.767602E-4   -3.000025E-5   1.792879E-4   -9.633516E+0   -9.632616E+0   
1.269260E+4   2.067571E+1   2.067571E+1   6.180000E+2   6.180000E+2   9.000000E-4   6.190000E+2   6.190000E+2   1.295764E-1   8.325547E-2   1.841373E-4   -3.964409E-5   1.841379E-4   -3.964120E-5   1.883565E-4   -1.215011E+1   -1.214921E+1   
1.272009E+4   2.068331E+1   2.068331E+1   6.280000E+2   6.280000E+2   9.000000E-4   6.290000E+2   6.290000E+2   1.328120E-1   8.128891E-2   1.856657E-4   -3.630371E-5   1.856663E-4   -3.630080E-5   1.891817E-4   -1.106361E+1   -1.106271E+1   
1.274707E+4   2.066171E+1   2.066171E+1   6.390000E+2   6.390000E+2   9.000000E-4   6.390000E+2   6.390000E+2   1.335487E-1   8.082392E-2   1.865143E-4   -3.555901E-5   1.865148E-4   -3.555608E-5   1.898737E-4   -1.079393E+1   -1.079303E+1   
1.277411E+4   2.066909E+1   2.066909E+1   6.480000E+2   6.480000E+2   9.000000E-4   6.490000E+2   6.490000E+2   1.328796E-1   8.446180E-2   1.892716E-4   -3.828795E-5   1.892722E-4   -3.828497E-5   1.931054E-4   -1.143609E+1   -1.143519E+1   
1.280107E+4   2.066601E+1   2.066601E+1   6.580000E+2   6.580000E+2   9.000000E-4   6.590000E+2   6.590000E+2   1.341743E-1   8.252814E-2   1.894749E-4   -3.626333E-5   1.894755E-4   -3.626036E-5   1.929139E-4   -1.083474E+1   -1.083384E+1   
1.282815E+4   2.067141E+1   2.067141E+1   6.680000E+2   6.680000E+2   9.000000E-4   6.690000E+2   6.690000E+2   1.349498E-1   8.381093E-2   1.915795E-4   -3.657281E-5   1.915801E-4   -3.656980E-5   1.950392E-4   -1.080781E+1   -1.080691E+1   
1.285525E+4   2.065688E+1   2.065688E+1   6.780000E+2   6.780000E+2   9.000000E-4   6.790000E+2   6.790000E+2   1.361686E-1   8.665806E-2   1.950922E-4   -3.755308E-5   1.950928E-4   -3.755001E-5   1.986736E-4   -1.089554E+1   -1.089464E+1   
1.288227E+4   2.064871E+1   2.064871E+1   6.880000E+2   6.880000E+2   9.000000E-4   6.890000E+2   6.890000E+2   1.368029E-1   8.497091E-2   1.950101E-4   -3.612148E-5   1.950107E-4   -3.611842E-5   1.983273E-4   -1.049389E+1   -1.049299E+1   
1.290932E+4   2.064050E+1   2.064050E+1   6.980000E+2   6.980000E+2   9.000000E-4   6.990000E+2   6.990000E+2   1.381872E-1   8.614249E-2   1.974594E-4   -3.595592E-5   1.974600E-4   -3.595282E-5   2.007064E-4   -1.032007E+1   -1.031917E+1   
1.293628E+4   2.065261E+1   2.065261E+1   7.080000E+2   7.080000E+2   9.000000E-4   7.090000E+2   7.090000E+2   1.382557E-1   8.823856E-2   1.996449E-4   -3.723979E-5   1.996455E-4   -3.723665E-5   2.030884E-4   -1.056596E+1   -1.056506E+1   
1.296331E+4   2.065869E+1   2.065869E+1   7.180000E+2   7.180000E+2   9.000000E-4   7.190000E+2   7.190000E+2   1.382856E-1   8.940526E-2   2.011499E-4   -3.797517E-5   2.011505E-4   -3.797201E-5   2.047032E-4   -1.069106E+1   -1.069016E+1   
1.299077E+4   2.064919E+1   2.064919E+1   7.280000E+2   7.280000E+2   9.000000E-4   7.280000E+2   7.280000E+2   1.398481E-1   8.929984E-2   2.027586E-4   -3.689811E-5   2.027592E-4   -3.689492E-5   2.060886E-4   -1.031385E+1   -1.031295E+1   
1.301818E+4   2.064300E+1   2.064300E+1   7.380000E+2   7.380000E+2   9.000000E-4   7.390000E+2   7.390000E+2   1.398432E-1   8.971240E-2   2.037755E-4   -3.719409E-5   2.037761E-4   -3.719089E-5   2.071421E-4   -1.034404E+1   -1.034314E+1   
1.304564E+4   2.063979E+1   2.063979E+1   7.480000E+2   7.480000E+2   9.000000E-4   7.490000E+2   7.490000E+2   1.402241E-1   9.048998E-2   2.052507E-4   -3.745476E-5   2.052513E-4   -3.745154E-5   2.086401E-4   -1.034172E+1   -1.034082E+1   
1.307312E+4   2.063769E+1   2.063769E+1   7.580000E+2   7.580000E+2   9.000000E-4   7.590000E+2   7.590000E+2   1.412662E-1   9.147052E-2   2.073279E-4   -3.739952E-5   2.073285E-4   -3.739627E-5   2.106741E-4   -1.022552E+1   -1.022462E+1   
1.310060E+4   2.064721E+1   2.064721E+1   7.680000E+2   7.680000E+2   9.000000E-4   7.690000E+2   7.690000E+2   1.423887E-1   9.142326E-2   2.087382E-4   -3.665549E-5   2.087388E-4   -3.665221E-5   2.119322E-4   -9.959879E+0   -9.958979E+0   
1.312808E+4   2.064681E+1   2.064681E+1   7.780000E+2   7.780000E+2   9.000000E-4   7.790000E+2   7.790000E+2   1.413292E-1   9.381274E-2   2.103465E-4   -3.887353E-5   2.103471E-4   -3.887022E-5   2.139084E-4   -1.047053E+1   -1.046963E+1   
1.315534E+4   2.066561E+1   2.066561E+1   7.880000E+2   7.880000E+2   9.000000E-4   7.890000E+2   7.890000E+2   1.438594E-1   9.520066E-2   2.137440E-4   -3.807680E-5   2.137446E-4   -3.807344E-5   2.171090E-4   -1.010083E+1   -1.009993E+1   
1.318228E+4   2.065551E+1   2.065551E+1   7.980000E+2   7.980000E+2   9.000000E-4   7.990000E+2   7.990000E+2   1.445021E-1   9.399039E-2   2.140030E-4   -3.693438E-5   2.140036E-4   -3.693102E-5   2.171668E-4   -9.792107E+0   -9.791207E+0   
1.320933E+4   2.067501E+1   2.067501E+1   8.080000E+2   8.080000E+2   9.000000E-4   8.090000E+2   8.090000E+2   1.445475E-1   9.594048E-2   2.160698E-4   -3.814349E-5   2.160704E-4   -3.814009E-5   2.194107E-4   -1.001146E+1   -1.001056E+1   
1.323638E+4   2.065399E+1   2.065399E+1   8.180000E+2   8.180000E+2   9.000000E-4   8.190000E+2   8.190000E+2   1.448147E-1   9.705933E-2   2.177060E-4   -3.869089E-5   2.177066E-4   -3.868747E-5   2.211173E-4   -1.007743E+1   -1.007653E+1   
1.326337E+4   2.065911E+1   2.065911E+1   8.280000E+2   8.280000E+2   9.000000E-4   8.290000E+2   8.290000E+2   1.475564E-1   9.756119E-2   2.206273E-4   -3.720549E-5   2.206279E-4   -3.720202E-5   2.237424E-4   -9.572018E+0   -9.571118E+0   
1.329087E+4   2.065630E+1   2.065630E+1   8.380000E+2   8.380000E+2   9.000000E-4   8.390000E+2   8.390000E+2   1.462297E-1   9.746397E-2   2.203011E-4   -3.806524E-5   2.203017E-4   -3.806178E-5   2.235655E-4   -9.803192E+0   -9.802292E+0   
1.331788E+4   2.066900E+1   2.066900E+1   8.480000E+2   8.480000E+2   9.000000E-4   8.490000E+2   8.490000E+2   1.470015E-1   9.778179E-2   2.217245E-4   -3.778088E-5   2.217251E-4   -3.777740E-5   2.249203E-4   -9.670075E+0   -9.669175E+0   
1.334532E+4   2.065789E+1   2.065789E+1   8.580000E+2   8.580000E+2   9.000000E-4   8.590000E+2   8.590000E+2   1.473208E-1   9.879159E-2   2.233203E-4   -3.822611E-5   2.233209E-4   -3.822260E-5   2.265682E-4   -9.713281E+0   -9.712381E+0   
1.337228E+4   2.067440E+1   2.067440E+1   8.680000E+2   8.680000E+2   9.000000E-4   8.690000E+2   8.690000E+2   1.451715E-1   9.780465E-2   2.217969E-4   -3.908515E-5   2.217975E-4   -3.908166E-5   2.252143E-4   -9.994081E+0   -9.993181E+0   
1.339982E+4   2.066580E+1   2.066580E+1   8.780000E+2   8.780000E+2   9.000000E-4   8.790000E+2   8.790000E+2   1.445094E-1   9.681680E-2   2.213060E-4   -3.895099E-5   2.213066E-4   -3.894751E-5   2.247076E-4   -9.982115E+0   -9.981215E+0   
1.342682E+4   2.067001E+1   2.067001E+1   8.880000E+2   8.880000E+2   9.000000E-4   8.890000E+2   8.890000E+2   1.455798E-1   9.852863E-2   2.239172E-4   -3.932874E-5   2.239178E-4   -3.932523E-5   2.273448E-4   -9.961804E+0   -9.960904E+0   
1.345388E+4   2.068401E+1   2.068401E+1   8.980000E+2   8.980000E+2   9.000000E-4   8.990000E+2   8.990000E+2   1.461212E-1   9.996285E-2   2.259657E-4   -3.988800E-5   2.259663E-4   -3.988445E-5   2.294593E-4   -1.001086E+1   -1.000996E+1   
1.348090E+4   2.066760E+1   2.066760E+1   9.080000E+2   9.080000E+2   9.000000E-4   9.090000E+2   9.090000E+2   1.451118E-1   1.007064E-1   2.264511E-4   -4.105554E-5   2.264518E-4   -4.105199E-5   2.301427E-4   -1.027609E+1   -1.027519E+1   
1.350834E+4   2.066851E+1   2.066851E+1   9.180000E+2   9.180000E+2   9.000000E-4   9.190000E+2   9.190000E+2   1.468123E-1   1.008480E-1   2.283958E-4   -4.004247E-5   2.283965E-4   -4.003888E-5   2.318794E-4   -9.944062E+0   -9.943162E+0   
1.353535E+4   2.066879E+1   2.066879E+1   9.280000E+2   9.280000E+2   9.000000E-4   9.290000E+2   9.290000E+2   1.468595E-1   1.015525E-1   2.295878E-4   -4.048064E-5   2.295884E-4   -4.047704E-5   2.331292E-4   -9.999545E+0   -9.998645E+0   
1.356285E+4   2.066281E+1   2.066281E+1   9.380000E+2   9.380000E+2   9.000000E-4   9.390000E+2   9.390000E+2   1.485012E-1   1.009166E-1   2.309448E-4   -3.902631E-5   2.309454E-4   -3.902268E-5   2.342190E-4   -9.591538E+0   -9.590638E+0   
1.358989E+4   2.066381E+1   2.066381E+1   9.480000E+2   9.480000E+2   9.000000E-4   9.490000E+2   9.490000E+2   1.474433E-1   1.015763E-1   2.313376E-4   -4.017442E-5   2.313383E-4   -4.017078E-5   2.348001E-4   -9.851811E+0   -9.850911E+0   
1.361695E+4   2.065341E+1   2.065341E+1   9.590000E+2   9.590000E+2   9.000000E-4   9.590000E+2   9.590000E+2   1.499854E-1   1.019702E-1   2.340444E-4   -3.875555E-5   2.340450E-4   -3.875188E-5   2.372315E-4   -9.402324E+0   -9.401424E+0   
1.364450E+4   2.066091E+1   2.066091E+1   9.680000E+2   9.680000E+2   9.000000E-4   9.690000E+2   9.690000E+2   1.490104E-1   1.035361E-1   2.351321E-4   -4.040832E-5   2.351327E-4   -4.040463E-5   2.385790E-4   -9.751241E+0   -9.750341E+0   
1.367148E+4   2.066851E+1   2.066851E+1   9.780000E+2   9.780000E+2   9.000000E-4   9.790000E+2   9.790000E+2   1.496040E-1   1.035230E-1   2.361990E-4   -4.003843E-5   2.361996E-4   -4.003472E-5   2.395684E-4   -9.620838E+0   -9.619938E+0   
1.369902E+4   2.066311E+1   2.066311E+1   9.880000E+2   9.880000E+2   9.000000E-4   9.890000E+2   9.890000E+2   1.499519E-1   1.054826E-1   2.384825E-4   -4.105144E-5   2.384832E-4   -4.104770E-5   2.419899E-4   -9.766954E+0   -9.766054E+0   
1.372603E+4   2.066250E+1   2.066250E+1   9.980000E+2   9.980000E+2   9.000000E-4   9.990000E+2   9.990000E+2   1.505613E-1   1.058522E-1   2.398295E-4   -4.090748E-5   2.398302E-4   -4.090371E-5   2.432933E-4   -9.679726E+0   -9.678826E+0   
1.375367E+4   2.066320E+1   2.066320E+1   1.008000E+3   1.008000E+3   9.000000E-4   1.009000E+3   1.009000E+3   1.518563E-1   1.055179E-1   2.411578E-4   -3.987100E-5   2.411585E-4   -3.986721E-5   2.444316E-4   -9.387878E+0   -9.386978E+0   
1.378109E+4   2.066091E+1   2.066091E+1   1.018000E+3   1.018000E+3   9.000000E-4   1.019000E+3   1.019000E+3   1.524909E-1   1.071478E-1   2.434087E-4   -4.048892E-5   2.434093E-4   -4.048509E-5   2.467532E-4   -9.444182E+0   -9.443282E+0   
1.380878E+4   2.066119E+1   2.066119E+1   1.028000E+3   1.028000E+3   9.000000E-4   1.029000E+3   1.029000E+3   1.537012E-1   1.076688E-1   2.452796E-4   -4.003748E-5   2.452803E-4   -4.003362E-5   2.485259E-4   -9.270741E+0   -9.269841E+0   
1.383618E+4   2.066790E+1   2.066790E+1   1.039000E+3   1.039000E+3   9.000000E-4   1.039000E+3   1.039000E+3   1.552043E-1   1.081530E-1   2.473281E-4   -3.936783E-5   2.473287E-4   -3.936395E-5   2.504416E-4   -9.044043E+0   -9.043143E+0   
1.386391E+4   2.066741E+1   2.066741E+1   1.048000E+3   1.048000E+3   9.000000E-4   1.049000E+3   1.049000E+3   1.554764E-1   1.085521E-1   2.484615E-4   -3.946724E-5   2.484622E-4   -3.946333E-5   2.515766E-4   -9.025822E+0   -9.024922E+0   
1.389137E+4   2.068731E+1   2.068731E+1   1.058000E+3   1.058000E+3   9.000000E-4   1.059000E+3   1.059000E+3   1.575173E-1   1.062940E-1   2.489550E-4   -3.674409E-5   2.489556E-4   -3.674018E-5   2.516520E-4   -8.395858E+0   -8.394958E+0   
1.391907E+4   2.068920E+1   2.068920E+1   1.068000E+3   1.068000E+3   9.000000E-4   1.069000E+3   1.069000E+3   1.508313E-1   1.125632E-1   2.493831E-4   -4.511488E-5   2.493838E-4   -4.511097E-5   2.534310E-4   -1.025424E+1   -1.025334E+1   
1.394647E+4   2.067809E+1   2.067809E+1   1.079000E+3   1.079000E+3   9.000000E-4   1.079000E+3   1.079000E+3   1.557558E-1   1.131650E-1   2.538910E-4   -4.223432E-5   2.538916E-4   -4.223033E-5   2.573798E-4   -9.444571E+0   -9.443671E+0   
1.397421E+4   2.067599E+1   2.067599E+1   1.088000E+3   1.088000E+3   9.000000E-4   1.089000E+3   1.089000E+3   1.589789E-1   1.138463E-1   2.572729E-4   -4.053850E-5   2.572735E-4   -4.053446E-5   2.604471E-4   -8.954475E+0   -8.953575E+0   
1.400163E+4   2.066689E+1   2.066689E+1   1.098000E+3   1.098000E+3   9.000000E-4   1.099000E+3   1.099000E+3   1.597138E-1   1.117210E-1   2.569526E-4   -3.876906E-5   2.569532E-4   -3.876502E-5   2.598609E-4   -8.580081E+0   -8.579181E+0   
1.402912E+4   2.068151E+1   2.068151E+1   1.108000E+3   1.108000E+3   9.000000E-4   1.109000E+3   1.109000E+3   1.584146E-1   1.125870E-1   2.573228E-4   -4.020568E-5   2.573234E-4   -4.020164E-5   2.604448E-4   -8.880441E+0   -8.879541E+0   
1.405683E+4   2.068130E+1   2.068130E+1   1.119000E+3   1.119000E+3   9.000000E-4   1.119000E+3   1.119000E+3   1.620570E-1   1.172738E-1   2.638129E-4   -4.070523E-5   2.638135E-4   -4.070109E-5   2.669348E-4   -8.771329E+0   -8.770429E+0   
1.408433E+4   2.067300E+1   2.067300E+1   1.128000E+3   1.128000E+3   9.000000E-4   1.129000E+3   1.129000E+3   1.581334E-1   1.188169E-1   2.628362E-4   -4.431181E-5   2.628369E-4   -4.430768E-5   2.665453E-4   -9.569563E+0   -9.568663E+0   
1.411205E+4   2.068121E+1   2.068121E+1   1.138000E+3   1.138000E+3   9.000000E-4   1.139000E+3   1.139000E+3   1.599302E-1   1.072237E-1   2.565951E-4   -3.598302E-5   2.565957E-4   -3.597899E-5   2.591059E-4   -7.982685E+0   -7.981785E+0   
1.413954E+4   2.068551E+1   2.068551E+1   1.148000E+3   1.148000E+3   9.000000E-4   1.149000E+3   1.149000E+3   1.620052E-1   1.179454E-1   2.662405E-4   -4.125788E-5   2.662412E-4   -4.125370E-5   2.694183E-4   -8.808759E+0   -8.807859E+0   
1.416723E+4   2.068139E+1   2.068139E+1   1.159000E+3   1.159000E+3   9.000000E-4   1.159000E+3   1.159000E+3   1.605064E-1   1.176060E-1   2.656244E-4   -4.208285E-5   2.656251E-4   -4.207868E-5   2.689373E-4   -9.002541E+0   -9.001641E+0   
1.419472E+4   2.067001E+1   2.067001E+1   1.169000E+3   1.169000E+3   9.000000E-4   1.169000E+3   1.169000E+3   1.611566E-1   1.157979E-1   2.654683E-4   -4.056595E-5   2.654690E-4   -4.056178E-5   2.685499E-4   -8.688102E+0   -8.687202E+0   
1.422240E+4   2.067681E+1   2.067681E+1   1.178000E+3   1.178000E+3   9.000000E-4   1.179000E+3   1.179000E+3   1.628270E-1   1.157302E-1   2.672449E-4   -3.944367E-5   2.672455E-4   -3.943947E-5   2.701400E-4   -8.395884E+0   -8.394984E+0   
1.424958E+4   2.067550E+1   2.067550E+1   1.188000E+3   1.188000E+3   9.000000E-4   1.189000E+3   1.189000E+3   1.625098E-1   1.160593E-1   2.679197E-4   -3.989308E-5   2.679203E-4   -3.988887E-5   2.708735E-4   -8.469082E+0   -8.468182E+0   
1.427727E+4   2.068130E+1   2.068130E+1   1.199000E+3   1.199000E+3   9.000000E-4   1.199000E+3   1.199000E+3   1.619854E-1   1.197715E-1   2.708298E-4   -4.257133E-5   2.708305E-4   -4.256707E-5   2.741553E-4   -8.933142E+0   -8.932242E+0   
1.430466E+4   2.067199E+1   2.067199E+1   1.209000E+3   1.209000E+3   9.000000E-4   1.209000E+3   1.209000E+3   1.620381E-1   1.185734E-1   2.706877E-4   -4.183019E-5   2.706883E-4   -4.182594E-5   2.739007E-4   -8.784605E+0   -8.783705E+0   
1.433234E+4   2.067251E+1   2.067251E+1   1.219000E+3   1.219000E+3   9.000000E-4   1.219000E+3   1.219000E+3   1.628818E-1   1.219336E-1   2.743006E-4   -4.337785E-5   2.743013E-4   -4.337354E-5   2.777093E-4   -8.986326E+0   -8.985426E+0   
1.435980E+4   2.066729E+1   2.066729E+1   1.228000E+3   1.228000E+3   9.000000E-4   1.229000E+3   1.229000E+3   1.637038E-1   1.215896E-1   2.752935E-4   -4.265098E-5   2.752942E-4   -4.264665E-5   2.785779E-4   -8.806766E+0   -8.805866E+0   
1.438751E+4   2.068020E+1   2.068020E+1   1.239000E+3   1.239000E+3   9.000000E-4   1.239000E+3   1.239000E+3   1.650034E-1   1.194232E-1   2.753365E-4   -4.047926E-5   2.753372E-4   -4.047494E-5   2.782962E-4   -8.363563E+0   -8.362663E+0   
1.441493E+4   2.067321E+1   2.067321E+1   1.248000E+3   1.248000E+3   9.000000E-4   1.249000E+3   1.249000E+3   1.666366E-1   1.215479E-1   2.786290E-4   -4.073649E-5   2.786297E-4   -4.073212E-5   2.815912E-4   -8.317902E+0   -8.317002E+0   
1.444262E+4   2.066390E+1   2.066390E+1   1.259000E+3   1.259000E+3   9.000000E-4   1.259000E+3   1.259000E+3   1.664035E-1   1.216021E-1   2.791690E-4   -4.095996E-5   2.791696E-4   -4.095557E-5   2.821578E-4   -8.346940E+0   -8.346040E+0   
1.447010E+4   2.065609E+1   2.065609E+1   1.268000E+3   1.268000E+3   9.000000E-4   1.269000E+3   1.269000E+3   1.666866E-1   1.260586E-1   2.831635E-4   -4.355927E-5   2.831642E-4   -4.355482E-5   2.864943E-4   -8.745302E+0   -8.744402E+0   
1.449729E+4   2.066790E+1   2.066790E+1   1.279000E+3   1.279000E+3   9.000000E-4   1.280000E+3   1.280000E+3   1.674998E-1   1.245370E-1   2.833885E-4   -4.211398E-5   2.833891E-4   -4.210953E-5   2.865006E-4   -8.452787E+0   -8.451887E+0   
1.452494E+4   2.065750E+1   2.065750E+1   1.288000E+3   1.288000E+3   9.000000E-4   1.289000E+3   1.289000E+3   1.657674E-1   1.236725E-1   2.821745E-4   -4.276705E-5   2.821751E-4   -4.276262E-5   2.853970E-4   -8.618297E+0   -8.617397E+0   
1.455233E+4   2.066940E+1   2.066940E+1   1.298000E+3   1.298000E+3   9.000000E-4   1.299000E+3   1.299000E+3   1.662241E-1   1.168448E-1   2.783539E-4   -3.827746E-5   2.783545E-4   -3.827309E-5   2.809734E-4   -7.829844E+0   -7.828944E+0   
1.458003E+4   2.065530E+1   2.065530E+1   1.308000E+3   1.308000E+3   9.000000E-4   1.309000E+3   1.309000E+3   1.670955E-1   1.254468E-1   2.856724E-4   -4.304570E-5   2.856731E-4   -4.304122E-5   2.888973E-4   -8.568980E+0   -8.568080E+0   
1.460752E+4   2.064669E+1   2.064669E+1   1.319000E+3   1.319000E+3   9.000000E-4   1.319000E+3   1.319000E+3   1.682705E-1   1.255501E-1   2.872250E-4   -4.235972E-5   2.872257E-4   -4.235521E-5   2.903318E-4   -8.389462E+0   -8.388562E+0   
1.463522E+4   2.064221E+1   2.064221E+1   1.329000E+3   1.329000E+3   9.000000E-4   1.329000E+3   1.329000E+3   1.691894E-1   1.288143E-1   2.908228E-4   -4.379785E-5   2.908235E-4   -4.379329E-5   2.941023E-4   -8.564373E+0   -8.563473E+0   
1.466258E+4   2.064150E+1   2.064150E+1   1.338000E+3   1.338000E+3   9.000000E-4   1.339000E+3   1.339000E+3   1.696498E-1   1.272634E-1   2.907157E-4   -4.256655E-5   2.907163E-4   -4.256198E-5   2.938154E-4   -8.330049E+0   -8.329149E+0   
1.469032E+4   2.066430E+1   2.066430E+1   1.348000E+3   1.348000E+3   9.000000E-4   1.349000E+3   1.349000E+3   1.698146E-1   1.269081E-1   2.912441E-4   -4.227137E-5   2.912447E-4   -4.226680E-5   2.942957E-4   -8.258283E+0   -8.257383E+0   
1.471777E+4   2.065460E+1   2.065460E+1   1.359000E+3   1.359000E+3   9.000000E-4   1.359000E+3   1.359000E+3   1.674331E-1   1.294743E-1   2.920582E-4   -4.548100E-5   2.920589E-4   -4.547641E-5   2.955782E-4   -8.851339E+0   -8.850439E+0   
1.474552E+4   2.065429E+1   2.065429E+1   1.368000E+3   1.368000E+3   9.000000E-4   1.369000E+3   1.369000E+3   1.699646E-1   1.273030E-1   2.929535E-4   -4.248405E-5   2.929542E-4   -4.247945E-5   2.960180E-4   -8.251497E+0   -8.250597E+0   
1.477299E+4   2.064999E+1   2.064999E+1   1.378000E+3   1.378000E+3   9.000000E-4   1.379000E+3   1.379000E+3   1.705892E-1   1.287440E-1   2.950645E-4   -4.299198E-5   2.950652E-4   -4.298734E-5   2.981801E-4   -8.289870E+0   -8.288970E+0   
1.480063E+4   2.064889E+1   2.064889E+1   1.389000E+3   1.389000E+3   9.000000E-4   1.389000E+3   1.389000E+3   1.716614E-1   1.284380E-1   2.962580E-4   -4.212166E-5   2.962586E-4   -4.211700E-5   2.992374E-4   -8.092020E+0   -8.091120E+0   
1.482807E+4   2.066689E+1   2.066689E+1   1.399000E+3   1.399000E+3   9.000000E-4   1.400000E+3   1.400000E+3   1.718174E-1   1.276830E-1   2.965655E-4   -4.158875E-5   2.965662E-4   -4.158409E-5   2.994674E-4   -7.982793E+0   -7.981893E+0   
1.485531E+4   2.066680E+1   2.066680E+1   1.409000E+3   1.409000E+3   9.000000E-4   1.410000E+3   1.410000E+3   1.718655E-1   1.281620E-1   2.975996E-4   -4.188698E-5   2.976002E-4   -4.188231E-5   3.005329E-4   -8.011722E+0   -8.010822E+0   
1.488273E+4   2.066729E+1   2.066729E+1   1.419000E+3   1.419000E+3   9.000000E-4   1.419000E+3   1.419000E+3   1.721922E-1   1.303951E-1   2.999943E-4   -4.307984E-5   2.999950E-4   -4.307512E-5   3.030717E-4   -8.171931E+0   -8.171031E+0   
1.490996E+4   2.065420E+1   2.065420E+1   1.429000E+3   1.429000E+3   9.000000E-4   1.429000E+3   1.429000E+3   1.742992E-1   1.315694E-1   3.029476E-4   -4.243361E-5   3.029483E-4   -4.242885E-5   3.059050E-4   -7.973495E+0   -7.972595E+0   
1.493718E+4   2.066061E+1   2.066061E+1   1.439000E+3   1.439000E+3   9.000000E-4   1.440000E+3   1.440000E+3   1.765397E-1   1.337471E-1   3.067656E-4   -4.232172E-5   3.067663E-4   -4.231690E-5   3.096713E-4   -7.855002E+0   -7.854102E+0   
1.496460E+4   2.064779E+1   2.064779E+1   1.449000E+3   1.449000E+3   9.000000E-4   1.449000E+3   1.449000E+3   1.775065E-1   1.346950E-1   3.087013E-4   -4.229308E-5   3.087020E-4   -4.228823E-5   3.115850E-4   -7.801141E+0   -7.800241E+0   
1.499220E+4   2.067129E+1   2.067129E+1   1.459000E+3   1.459000E+3   9.000000E-4   1.460000E+3   1.460000E+3   1.790404E-1   1.357081E-1   3.112095E-4   -4.193317E-5   3.112101E-4   -4.192828E-5   3.140219E-4   -7.673962E+0   -7.673062E+0   
1.501943E+4   2.064419E+1   2.064419E+1   1.469000E+3   1.469000E+3   9.000000E-4   1.470000E+3   1.470000E+3   1.800340E-1   1.373032E-1   3.136852E-4   -4.229008E-5   3.136859E-4   -4.228515E-5   3.165231E-4   -7.678145E+0   -7.677245E+0   
1.504666E+4   2.063561E+1   2.063561E+1   1.479000E+3   1.479000E+3   9.000000E-4   1.480000E+3   1.480000E+3   1.817218E-1   1.389206E-1   3.166589E-4   -4.219737E-5   3.166596E-4   -4.219240E-5   3.194581E-4   -7.590409E+0   -7.589509E+0   
1.507388E+4   2.064099E+1   2.064099E+1   1.489000E+3   1.489000E+3   9.000000E-4   1.490000E+3   1.490000E+3   1.842415E-1   1.392759E-1   3.193229E-4   -4.076957E-5   3.193235E-4   -4.076456E-5   3.219150E-4   -7.275879E+0   -7.274979E+0   
1.510106E+4   2.063799E+1   2.063799E+1   1.499000E+3   1.499000E+3   9.000000E-4   1.499000E+3   1.499000E+3   1.845078E-1   1.402363E-1   3.207807E-4   -4.121624E-5   3.207813E-4   -4.121120E-5   3.234177E-4   -7.321664E+0   -7.320764E+0   
1.512822E+4   2.064761E+1   2.064761E+1   1.509000E+3   1.509000E+3   9.000000E-4   1.510000E+3   1.510000E+3   1.837780E-1   1.402634E-1   3.210229E-4   -4.175785E-5   3.210236E-4   -4.175281E-5   3.237274E-4   -7.411276E+0   -7.410376E+0   
1.515542E+4   2.064849E+1   2.064849E+1   1.519000E+3   1.519000E+3   9.000000E-4   1.520000E+3   1.520000E+3   1.842902E-1   1.412972E-1   3.227696E-4   -4.208922E-5   3.227702E-4   -4.208415E-5   3.255022E-4   -7.429460E+0   -7.428560E+0   
1.518266E+4   2.064370E+1   2.064370E+1   1.529000E+3   1.529000E+3   9.000000E-4   1.530000E+3   1.530000E+3   1.845513E-1   1.396089E-1   3.224274E-4   -4.090602E-5   3.224281E-4   -4.090096E-5   3.250119E-4   -7.230427E+0   -7.229527E+0   
1.520984E+4   2.063711E+1   2.063711E+1   1.539000E+3   1.539000E+3   9.000000E-4   1.540000E+3   1.540000E+3   1.850864E-1   1.414831E-1   3.247809E-4   -4.174141E-5   3.247816E-4   -4.173631E-5   3.274523E-4   -7.323607E+0   -7.322707E+0   
1.523703E+4   2.063070E+1   2.063070E+1   1.549000E+3   1.549000E+3   9.000000E-4   1.549000E+3   1.549000E+3   1.849332E-1   1.426580E-1   3.260981E-4   -4.260066E-5   3.260988E-4   -4.259553E-5   3.288690E-4   -7.442830E+0   -7.441930E+0   
1.526428E+4   2.063339E+1   2.063339E+1   1.559000E+3   1.559000E+3   9.000000E-4   1.559000E+3   1.559000E+3   1.857065E-1   1.413094E-1   3.263507E-4   -4.128551E-5   3.263514E-4   -4.128038E-5   3.289518E-4   -7.209992E+0   -7.209092E+0   
1.529142E+4   2.062829E+1   2.062829E+1   1.569000E+3   1.569000E+3   9.000000E-4   1.570000E+3   1.570000E+3   1.847168E-1   1.422479E-1   3.270534E-4   -4.256379E-5   3.270540E-4   -4.255865E-5   3.298114E-4   -7.414984E+0   -7.414084E+0   
1.531862E+4   2.063671E+1   2.063671E+1   1.579000E+3   1.579000E+3   9.000000E-4   1.580000E+3   1.580000E+3   1.845068E-1   1.411677E-1   3.268116E-4   -4.207084E-5   3.268123E-4   -4.206570E-5   3.295084E-4   -7.335409E+0   -7.334509E+0   
1.534589E+4   2.062179E+1   2.062179E+1   1.589000E+3   1.589000E+3   9.000000E-4   1.590000E+3   1.590000E+3   1.851050E-1   1.424542E-1   3.287956E-4   -4.250091E-5   3.287963E-4   -4.249574E-5   3.315311E-4   -7.365348E+0   -7.364448E+0   
1.537306E+4   2.062591E+1   2.062591E+1   1.599000E+3   1.599000E+3   9.000000E-4   1.600000E+3   1.600000E+3   1.854103E-1   1.434076E-1   3.303420E-4   -4.292065E-5   3.303427E-4   -4.291546E-5   3.331186E-4   -7.402851E+0   -7.401951E+0   
1.540021E+4   2.062600E+1   2.062600E+1   1.609000E+3   1.609000E+3   9.000000E-4   1.610000E+3   1.610000E+3   1.867964E-1   1.419898E-1   3.309716E-4   -4.115380E-5   3.309722E-4   -4.114860E-5   3.335203E-4   -7.087915E+0   -7.087015E+0   
1.542744E+4   2.062011E+1   2.062011E+1   1.619000E+3   1.619000E+3   9.000000E-4   1.619000E+3   1.619000E+3   1.828885E-1   1.467547E-1   3.322053E-4   -4.673737E-5   3.322060E-4   -4.673215E-5   3.354768E-4   -8.008282E+0   -8.007382E+0   
1.545467E+4   2.062621E+1   2.062621E+1   1.629000E+3   1.629000E+3   9.000000E-4   1.630000E+3   1.630000E+3   1.861553E-1   1.420544E-1   3.318992E-4   -4.169033E-5   3.318999E-4   -4.168512E-5   3.345073E-4   -7.159507E+0   -7.158607E+0   
1.548189E+4   2.062960E+1   2.062960E+1   1.639000E+3   1.639000E+3   9.000000E-4   1.639000E+3   1.639000E+3   1.847908E-1   1.354619E-1   3.269125E-4   -3.855823E-5   3.269131E-4   -3.855309E-5   3.291785E-4   -6.726766E+0   -6.725866E+0   
1.550906E+4   2.063351E+1   2.063351E+1   1.649000E+3   1.649000E+3   9.000000E-4   1.650000E+3   1.650000E+3   1.923545E-1   1.468653E-1   3.409165E-4   -4.059436E-5   3.409171E-4   -4.058900E-5   3.433248E-4   -6.790477E+0   -6.789577E+0   
1.553627E+4   2.064611E+1   2.064611E+1   1.659000E+3   1.659000E+3   9.000000E-4   1.660000E+3   1.660000E+3   2.008115E-1   1.388517E-1   3.418194E-4   -3.003240E-5   3.418198E-4   -3.002704E-5   3.431362E-4   -5.021139E+0   -5.020239E+0   
1.556340E+4   2.062261E+1   2.062261E+1   1.669000E+3   1.669000E+3   9.000000E-4   1.670000E+3   1.670000E+3   1.893961E-1   1.458028E-1   3.394417E-4   -4.198106E-5   3.394423E-4   -4.197573E-5   3.420279E-4   -7.050358E+0   -7.049458E+0   
1.559059E+4   2.062191E+1   2.062191E+1   1.679000E+3   1.679000E+3   9.000000E-4   1.680000E+3   1.680000E+3   1.887413E-1   1.575858E-1   3.479371E-4   -4.973371E-5   3.479378E-4   -4.972824E-5   3.514735E-4   -8.134687E+0   -8.133787E+0   
1.561783E+4   2.062771E+1   2.062771E+1   1.689000E+3   1.689000E+3   9.000000E-4   1.689000E+3   1.689000E+3   1.895372E-1   1.460935E-1   3.410053E-4   -4.213180E-5   3.410060E-4   -4.212645E-5   3.435982E-4   -7.043300E+0   -7.042400E+0   
1.564507E+4   2.063540E+1   2.063540E+1   1.699000E+3   1.699000E+3   9.000000E-4   1.699000E+3   1.699000E+3   1.956201E-1   1.652773E-1   3.593859E-4   -4.996073E-5   3.593867E-4   -4.995509E-5   3.628420E-4   -7.914362E+0   -7.913462E+0   
1.567221E+4   2.062161E+1   2.062161E+1   1.709000E+3   1.709000E+3   9.000000E-4   1.710000E+3   1.710000E+3   1.897807E-1   1.549544E-1   3.487999E-4   -4.751704E-5   3.488006E-4   -4.751156E-5   3.520216E-4   -7.757654E+0   -7.756754E+0   
1.569940E+4   2.063790E+1   2.063790E+1   1.719000E+3   1.719000E+3   9.000000E-4   1.720000E+3   1.720000E+3   1.908483E-1   1.456102E-1   3.436339E-4   -4.106465E-5   3.436346E-4   -4.105925E-5   3.460789E-4   -6.814595E+0   -6.813695E+0   
1.572711E+4   2.061700E+1   2.061700E+1   1.729000E+3   1.729000E+3   9.000000E-4   1.729000E+3   1.729000E+3   1.913712E-1   1.503130E-1   3.479018E-4   -4.365260E-5   3.479025E-4   -4.364713E-5   3.506297E-4   -7.151750E+0   -7.150850E+0   
1.575422E+4   2.062811E+1   2.062811E+1   1.739000E+3   1.739000E+3   9.000000E-4   1.740000E+3   1.740000E+3   1.921577E-1   1.557869E-1   3.530279E-4   -4.654804E-5   3.530286E-4   -4.654250E-5   3.560834E-4   -7.511334E+0   -7.510434E+0   
1.578141E+4   2.062829E+1   2.062829E+1   1.749000E+3   1.749000E+3   9.000000E-4   1.750000E+3   1.750000E+3   1.908091E-1   1.510092E-1   3.493948E-4   -4.453021E-5   3.493955E-4   -4.452472E-5   3.522211E-4   -7.263163E+0   -7.262263E+0   
1.580860E+4   2.063210E+1   2.063210E+1   1.759000E+3   1.759000E+3   9.000000E-4   1.760000E+3   1.760000E+3   1.923356E-1   1.495741E-1   3.501098E-4   -4.265889E-5   3.501104E-4   -4.265339E-5   3.526991E-4   -6.946924E+0   -6.946024E+0   
1.583578E+4   2.063641E+1   2.063641E+1   1.769000E+3   1.769000E+3   9.000000E-4   1.770000E+3   1.770000E+3   1.913060E-1   1.506384E-1   3.508068E-4   -4.403813E-5   3.508075E-4   -4.403262E-5   3.535601E-4   -7.155131E+0   -7.154231E+0   
1.586293E+4   2.063821E+1   2.063821E+1   1.779000E+3   1.779000E+3   9.000000E-4   1.780000E+3   1.780000E+3   1.932896E-1   1.445730E-1   3.485830E-4   -3.900056E-5   3.485836E-4   -3.899509E-5   3.507580E-4   -6.383882E+0   -6.382982E+0   
1.589017E+4   2.062661E+1   2.062661E+1   1.789000E+3   1.789000E+3   9.000000E-4   1.790000E+3   1.790000E+3   1.909294E-1   1.601389E-1   3.585541E-4   -5.022899E-5   3.585548E-4   -5.022336E-5   3.620552E-4   -7.974535E+0   -7.973635E+0   
1.591731E+4   2.063320E+1   2.063320E+1   1.799000E+3   1.799000E+3   9.000000E-4   1.800000E+3   1.800000E+3   1.880926E-1   1.543183E-1   3.531537E-4   -4.855990E-5   3.531545E-4   -4.855435E-5   3.564767E-4   -7.829277E+0   -7.828377E+0   
1.594451E+4   2.062609E+1   2.062609E+1   1.809000E+3   1.809000E+3   9.000000E-4   1.810000E+3   1.810000E+3   1.933158E-1   1.539867E-1   3.572128E-4   -4.490326E-5   3.572135E-4   -4.489765E-5   3.600240E-4   -7.164757E+0   -7.163857E+0   
1.597174E+4   2.062161E+1   2.062161E+1   1.819000E+3   1.819000E+3   9.000000E-4   1.820000E+3   1.820000E+3   1.928216E-1   1.484324E-1   3.536271E-4   -4.183520E-5   3.536278E-4   -4.182965E-5   3.560931E-4   -6.746913E+0   -6.746013E+0   
1.599897E+4   2.062499E+1   2.062499E+1   1.829000E+3   1.829000E+3   9.000000E-4   1.829000E+3   1.829000E+3   1.927464E-1   1.535333E-1   3.577595E-4   -4.506846E-5   3.577603E-4   -4.506284E-5   3.605871E-4   -7.179967E+0   -7.179067E+0   
1.602613E+4   2.062841E+1   2.062841E+1   1.839000E+3   1.839000E+3   9.000000E-4   1.840000E+3   1.840000E+3   1.916192E-1   1.512398E-1   3.560938E-4   -4.444131E-5   3.560945E-4   -4.443572E-5   3.588562E-4   -7.113862E+0   -7.112962E+0   
1.605328E+4   2.062380E+1   2.062380E+1   1.849000E+3   1.849000E+3   9.000000E-4   1.850000E+3   1.850000E+3   1.932217E-1   1.570380E-1   3.619483E-4   -4.698904E-5   3.619491E-4   -4.698335E-5   3.649857E-4   -7.396912E+0   -7.396012E+0   
1.608049E+4   2.061700E+1   2.061700E+1   1.859000E+3   1.859000E+3   9.000000E-4   1.860000E+3   1.860000E+3   1.951087E-1   1.509760E-1   3.596598E-4   -4.201798E-5   3.596605E-4   -4.201233E-5   3.621059E-4   -6.663489E+0   -6.662589E+0   
1.610769E+4   2.061389E+1   2.061389E+1   1.869000E+3   1.869000E+3   9.000000E-4   1.870000E+3   1.870000E+3   1.947669E-1   1.541823E-1   3.623410E-4   -4.426183E-5   3.623417E-4   -4.425614E-5   3.650344E-4   -6.964471E+0   -6.963571E+0   
1.613489E+4   2.061999E+1   2.061999E+1   1.879000E+3   1.879000E+3   9.000000E-4   1.880000E+3   1.880000E+3   1.939777E-1   1.547561E-1   3.628600E-4   -4.517750E-5   3.628607E-4   -4.517180E-5   3.656616E-4   -7.097029E+0   -7.096129E+0   
1.616211E+4   2.061971E+1   2.061971E+1   1.889000E+3   1.889000E+3   9.000000E-4   1.890000E+3   1.890000E+3   1.943573E-1   1.553737E-1   3.642219E-4   -4.534012E-5   3.642226E-4   -4.533440E-5   3.670331E-4   -7.095954E+0   -7.095054E+0   
1.618933E+4   2.062319E+1   2.062319E+1   1.899000E+3   1.899000E+3   9.000000E-4   1.900000E+3   1.900000E+3   1.943114E-1   1.553262E-1   3.648203E-4   -4.537580E-5   3.648210E-4   -4.537007E-5   3.676314E-4   -7.089951E+0   -7.089051E+0   
1.621655E+4   2.062850E+1   2.062850E+1   1.909000E+3   1.909000E+3   9.000000E-4   1.910000E+3   1.910000E+3   1.953278E-1   1.567126E-1   3.671652E-4   -4.558846E-5   3.671659E-4   -4.558269E-5   3.699845E-4   -7.077813E+0   -7.076913E+0   
1.624394E+4   2.063400E+1   2.063400E+1   1.919000E+3   1.919000E+3   9.000000E-4   1.920000E+3   1.920000E+3   1.966371E-1   1.548097E-1   3.674003E-4   -4.357309E-5   3.674010E-4   -4.356732E-5   3.699751E-4   -6.763595E+0   -6.762695E+0   
1.627109E+4   2.061440E+1   2.061440E+1   1.929000E+3   1.929000E+3   9.000000E-4   1.930000E+3   1.930000E+3   1.940478E-1   1.569591E-1   3.677769E-4   -4.666385E-5   3.677776E-4   -4.665807E-5   3.707254E-4   -7.231100E+0   -7.230200E+0   
1.629825E+4   2.061929E+1   2.061929E+1   1.939000E+3   1.939000E+3   9.000000E-4   1.940000E+3   1.940000E+3   1.980059E-1   1.572513E-1   3.713957E-4   -4.423700E-5   3.713964E-4   -4.423116E-5   3.740210E-4   -6.792507E+0   -6.791607E+0   
1.632548E+4   2.061669E+1   2.061669E+1   1.949000E+3   1.949000E+3   9.000000E-4   1.950000E+3   1.950000E+3   1.964942E-1   1.572732E-1   3.710248E-4   -4.529385E-5   3.710255E-4   -4.528803E-5   3.737793E-4   -6.960098E+0   -6.959198E+0   
1.635267E+4   2.062411E+1   2.062411E+1   1.959000E+3   1.959000E+3   9.000000E-4   1.960000E+3   1.960000E+3   1.951173E-1   1.585152E-1   3.716055E-4   -4.701472E-5   3.716062E-4   -4.700888E-5   3.745678E-4   -7.210628E+0   -7.209728E+0   
1.637988E+4   2.063491E+1   2.063491E+1   1.969000E+3   1.969000E+3   9.000000E-4   1.970000E+3   1.970000E+3   1.964659E-1   1.567854E-1   3.719896E-4   -4.508008E-5   3.719903E-4   -4.507423E-5   3.747112E-4   -6.909774E+0   -6.908874E+0   
1.640713E+4   2.062841E+1   2.062841E+1   1.979000E+3   1.979000E+3   9.000000E-4   1.980000E+3   1.980000E+3   1.968248E-1   1.590728E-1   3.745113E-4   -4.628833E-5   3.745121E-4   -4.628245E-5   3.773610E-4   -7.045831E+0   -7.044931E+0   
1.643429E+4   2.063448E+1   2.063448E+1   1.989000E+3   1.989000E+3   9.000000E-4   1.990000E+3   1.990000E+3   1.965506E-1   1.601484E-1   3.757410E-4   -4.717039E-5   3.757418E-4   -4.716449E-5   3.786903E-4   -7.155457E+0   -7.154557E+0   
1.646143E+4   2.062631E+1   2.062631E+1   1.999000E+3   1.999000E+3   9.000000E-4   2.000000E+3   2.000000E+3   1.964595E-1   1.579926E-1   3.748255E-4   -4.593342E-5   3.748262E-4   -4.592754E-5   3.776295E-4   -6.986543E+0   -6.985643E+0   
1.650165E+4   2.061929E+1   2.061929E+1   2.099000E+3   2.099000E+3   9.000000E-4   2.100000E+3   2.100000E+3   1.986129E-1   1.682787E-1   3.901929E-4   -5.119607E-5   3.901937E-4   -5.118994E-5   3.935372E-4   -7.474913E+0   -7.474013E+0   
1.652954E+4   2.061770E+1   2.061770E+1   2.199000E+3   2.199000E+3   9.000000E-4   2.200000E+3   2.200000E+3   2.089107E-1   1.562988E-1   3.955592E-4   -3.726380E-5   3.955597E-4   -3.725758E-5   3.973105E-4   -5.381688E+0   -5.380788E+0   
1.655766E+4   2.062509E+1   2.062509E+1   2.299000E+3   2.299000E+3   9.000000E-4   2.300000E+3   2.300000E+3   1.933694E-1   1.525815E-1   3.887867E-4   -4.568305E-5   3.887874E-4   -4.567694E-5   3.914614E-4   -6.701615E+0   -6.700715E+0   
1.658629E+4   2.063510E+1   2.063510E+1   2.399000E+3   2.399000E+3   9.000000E-4   2.399000E+3   2.399000E+3   1.876133E-1   1.629945E-1   3.986825E-4   -5.629978E-5   3.986833E-4   -5.629352E-5   4.026380E-4   -8.037853E+0   -8.036953E+0   
1.661492E+4   2.062991E+1   2.062991E+1   2.499000E+3   2.499000E+3   9.000000E-4   2.499000E+3   2.499000E+3   1.899458E-1   1.706986E-1   4.123584E-4   -5.984729E-5   4.123594E-4   -5.984082E-5   4.166787E-4   -8.257916E+0   -8.257016E+0   
1.664338E+4   2.061639E+1   2.061639E+1   2.598000E+3   2.598000E+3   9.000000E-4   2.599000E+3   2.599000E+3   1.782673E-1   1.485247E-1   3.952895E-4   -5.428339E-5   3.952904E-4   -5.427718E-5   3.989993E-4   -7.819272E+0   -7.818372E+0   
1.667224E+4   2.061749E+1   2.061749E+1   2.698000E+3   2.698000E+3   9.000000E-4   2.699000E+3   2.699000E+3   1.857900E-1   1.466276E-1   4.058189E-4   -4.843392E-5   4.058197E-4   -4.842755E-5   4.086989E-4   -6.805979E+0   -6.805079E+0   
1.670089E+4   2.062570E+1   2.062570E+1   2.799000E+3   2.799000E+3   9.000000E-4   2.799000E+3   2.799000E+3   1.806268E-1   1.423481E-1   4.058603E-4   -4.957917E-5   4.058611E-4   -4.957280E-5   4.088774E-4   -6.964643E+0   -6.963743E+0   
1.672923E+4   2.061611E+1   2.061611E+1   2.898000E+3   2.898000E+3   9.000000E-4   2.899000E+3   2.899000E+3   1.746028E-1   1.509672E-1   4.143747E-4   -5.926952E-5   4.143757E-4   -5.926301E-5   4.185921E-4   -8.140011E+0   -8.139111E+0   
1.675803E+4   2.061279E+1   2.061279E+1   2.999000E+3   2.999000E+3   9.000000E-4   3.000000E+3   3.000000E+3   1.706106E-1   1.334055E-1   4.059553E-4   -5.142906E-5   4.059561E-4   -5.142269E-5   4.092000E-4   -7.220141E+0   -7.219241E+0   
1.678666E+4   2.062869E+1   2.062869E+1   3.098000E+3   3.098000E+3   9.000000E-4   3.099000E+3   3.099000E+3   1.624324E-1   1.322465E-1   4.060303E-4   -5.651140E-5   4.060312E-4   -5.650502E-5   4.099441E-4   -7.923539E+0   -7.922639E+0   
1.681485E+4   2.063271E+1   2.063271E+1   3.199000E+3   3.199000E+3   9.000000E-4   3.199000E+3   3.199000E+3   1.704901E-1   1.116710E-1   4.037957E-4   -3.876272E-5   4.037963E-4   -3.875638E-5   4.056519E-4   -5.483357E+0   -5.482457E+0   
1.684374E+4   2.061810E+1   2.061810E+1   3.299000E+3   3.299000E+3   9.000000E-4   3.299000E+3   3.299000E+3   1.619294E-1   1.215147E-1   4.114091E-4   -5.090285E-5   4.114099E-4   -5.089639E-5   4.145462E-4   -7.053249E+0   -7.052349E+0   
1.687242E+4   2.062551E+1   2.062551E+1   3.399000E+3   3.399000E+3   9.000000E-4   3.399000E+3   3.399000E+3   1.572376E-1   1.147247E-1   4.100125E-4   -5.018221E-5   4.100133E-4   -5.017577E-5   4.130720E-4   -6.977835E+0   -6.976935E+0   
1.690107E+4   2.061379E+1   2.061379E+1   3.499000E+3   3.499000E+3   9.000000E-4   3.499000E+3   3.499000E+3   1.522731E-1   1.096018E-1   4.095988E-4   -5.067365E-5   4.095996E-4   -5.066722E-5   4.127215E-4   -7.052531E+0   -7.051631E+0   
1.692944E+4   2.061791E+1   2.061791E+1   3.599000E+3   3.599000E+3   9.000000E-4   3.600000E+3   3.600000E+3   1.465798E-1   1.043305E-1   4.086409E-4   -5.156325E-5   4.086417E-4   -5.155683E-5   4.118812E-4   -7.191706E+0   -7.190806E+0   
1.695738E+4   2.062869E+1   2.062869E+1   3.699000E+3   3.699000E+3   9.000000E-4   3.700000E+3   3.700000E+3   1.421885E-1   9.613366E-2   4.064636E-4   -4.977268E-5   4.064644E-4   -4.976629E-5   4.094997E-4   -6.981283E+0   -6.980383E+0   
1.698548E+4   2.063381E+1   2.063381E+1   3.799000E+3   3.799000E+3   9.000000E-4   3.800000E+3   3.800000E+3   1.371031E-1   9.330450E-2   4.075790E-4   -5.176225E-5   4.075798E-4   -5.175584E-5   4.108528E-4   -7.237777E+0   -7.236877E+0   
1.701411E+4   2.062170E+1   2.062170E+1   3.899000E+3   3.899000E+3   9.000000E-4   3.900000E+3   3.900000E+3   1.355335E-1   8.950061E-2   4.104513E-4   -5.080289E-5   4.104521E-4   -5.079644E-5   4.135834E-4   -7.055798E+0   -7.054898E+0   
1.704216E+4   2.061459E+1   2.061459E+1   3.999000E+3   3.999000E+3   9.000000E-4   4.000000E+3   4.000000E+3   1.302553E-1   8.699784E-2   4.116623E-4   -5.312286E-5   4.116631E-4   -5.311640E-5   4.150758E-4   -7.353084E+0   -7.352184E+0   
1.707030E+4   2.062670E+1   2.062670E+1   4.099000E+3   4.099000E+3   9.000000E-4   4.100000E+3   4.100000E+3   1.271604E-1   7.852342E-2   4.101904E-4   -5.029542E-5   4.101912E-4   -5.028898E-5   4.132624E-4   -6.990418E+0   -6.989518E+0   
1.709898E+4   2.063470E+1   2.063470E+1   4.199000E+3   4.199000E+3   9.000000E-4   4.199000E+3   4.199000E+3   1.212389E-1   7.311378E-2   4.088439E-4   -5.124502E-5   4.088447E-4   -5.123860E-5   4.120430E-4   -7.144269E+0   -7.143369E+0   
1.712762E+4   2.063110E+1   2.063110E+1   4.299000E+3   4.299000E+3   9.000000E-4   4.299000E+3   4.299000E+3   1.168515E-1   7.066491E-2   4.107117E-4   -5.300369E-5   4.107125E-4   -5.299724E-5   4.141177E-4   -7.353564E+0   -7.352664E+0   
1.715629E+4   2.064169E+1   2.064169E+1   4.399000E+3   4.399000E+3   9.000000E-4   4.399000E+3   4.399000E+3   1.141223E-1   6.423851E-2   4.109341E-4   -5.119776E-5   4.109349E-4   -5.119131E-5   4.141112E-4   -7.101814E+0   -7.100914E+0   
1.718522E+4   2.064581E+1   2.064581E+1   4.498000E+3   4.498000E+3   9.000000E-4   4.499000E+3   4.499000E+3   1.085768E-1   5.971190E-2   4.105361E-4   -5.244552E-5   4.105369E-4   -5.243907E-5   4.138725E-4   -7.280039E+0   -7.279139E+0   
1.721387E+4   2.064239E+1   2.064239E+1   4.599000E+3   4.599000E+3   9.000000E-4   4.599000E+3   4.599000E+3   1.041117E-1   5.494118E-2   4.107170E-4   -5.282132E-5   4.107179E-4   -5.281486E-5   4.140997E-4   -7.328443E+0   -7.327543E+0   
1.724231E+4   2.063329E+1   2.063329E+1   4.698000E+3   4.698000E+3   9.000000E-4   4.699000E+3   4.699000E+3   9.977181E-2   4.899770E-2   4.101602E-4   -5.238881E-5   4.101610E-4   -5.238237E-5   4.134924E-4   -7.278845E+0   -7.277945E+0   
1.727143E+4   2.063922E+1   2.063922E+1   4.798000E+3   4.798000E+3   9.000000E-4   4.799000E+3   4.799000E+3   9.578904E-2   4.611402E-2   4.120032E-4   -5.360875E-5   4.120041E-4   -5.360228E-5   4.154763E-4   -7.413522E+0   -7.412622E+0   
1.729981E+4   2.062579E+1   2.062579E+1   4.898000E+3   4.898000E+3   9.000000E-4   4.899000E+3   4.899000E+3   9.228256E-2   4.128665E-2   4.128102E-4   -5.330972E-5   4.128111E-4   -5.330324E-5   4.162382E-4   -7.358371E+0   -7.357471E+0   
1.732819E+4   2.061300E+1   2.061300E+1   4.998000E+3   4.998000E+3   9.000000E-4   4.999000E+3   4.999000E+3   8.786712E-2   3.612224E-2   4.127488E-4   -5.340908E-5   4.127496E-4   -5.340260E-5   4.161900E-4   -7.373020E+0   -7.372120E+0   
1.735729E+4   2.063448E+1   2.063448E+1   5.098000E+3   5.098000E+3   9.000000E-4   5.099000E+3   5.099000E+3   8.447308E-2   3.182992E-2   4.140102E-4   -5.336564E-5   4.140110E-4   -5.335914E-5   4.174354E-4   -7.344889E+0   -7.343989E+0   
1.738569E+4   2.063439E+1   2.063439E+1   5.198000E+3   5.198000E+3   9.000000E-4   5.199000E+3   5.199000E+3   7.696616E-2   2.825427E-2   4.129185E-4   -5.651010E-5   4.129193E-4   -5.650362E-5   4.167674E-4   -7.792823E+0   -7.791923E+0   
1.741408E+4   2.063549E+1   2.063549E+1   5.298000E+3   5.298000E+3   9.000000E-4   5.299000E+3   5.299000E+3   7.378840E-2   2.091770E-2   4.121892E-4   -5.444113E-5   4.121900E-4   -5.443466E-5   4.157689E-4   -7.523964E+0   -7.523064E+0   
1.744294E+4   2.062200E+1   2.062200E+1   5.398000E+3   5.398000E+3   9.000000E-4   5.399000E+3   5.399000E+3   7.035353E-2   1.525484E-2   4.124584E-4   -5.357802E-5   4.124592E-4   -5.357154E-5   4.159237E-4   -7.401234E+0   -7.400334E+0   
1.747162E+4   2.062811E+1   2.062811E+1   5.498000E+3   5.498000E+3   9.000000E-4   5.499000E+3   5.499000E+3   6.645641E-2   1.116606E-2   4.135134E-4   -5.399612E-5   4.135143E-4   -5.398962E-5   4.170239E-4   -7.439526E+0   -7.438626E+0   
1.749983E+4   2.064059E+1   2.064059E+1   5.599000E+3   5.599000E+3   9.000000E-4   5.599000E+3   5.599000E+3   6.185419E-2   4.852052E-3   4.125137E-4   -5.350976E-5   4.125146E-4   -5.350328E-5   4.159698E-4   -7.390928E+0   -7.390028E+0   
1.752894E+4   2.064611E+1   2.064611E+1   5.698000E+3   5.698000E+3   9.000000E-4   5.699000E+3   5.699000E+3   5.917193E-2   -1.858693E-4   4.137452E-4   -5.253051E-5   4.137460E-4   -5.252401E-5   4.170666E-4   -7.235755E+0   -7.234855E+0   
1.755738E+4   2.063922E+1   2.063922E+1   5.798000E+3   5.798000E+3   9.000000E-4   5.799000E+3   5.799000E+3   5.324551E-2   -3.905346E-3   4.136503E-4   -5.453123E-5   4.136511E-4   -5.452473E-5   4.172292E-4   -7.509957E+0   -7.509057E+0   
1.758572E+4   2.064111E+1   2.064111E+1   5.898000E+3   5.898000E+3   9.000000E-4   5.899000E+3   5.899000E+3   4.898611E-2   -8.675134E-3   4.139748E-4   -5.477030E-5   4.139756E-4   -5.476380E-5   4.175822E-4   -7.536660E+0   -7.535760E+0   
1.761466E+4   2.065371E+1   2.065371E+1   5.998000E+3   5.998000E+3   9.000000E-4   5.999000E+3   5.999000E+3   4.516547E-2   -1.211764E-2   4.155374E-4   -5.553671E-5   4.155383E-4   -5.553018E-5   4.192323E-4   -7.612487E+0   -7.611587E+0   
@@END Data.
@Time at end of measurement: 18:57:27
@Instrument  Changes:
@Emu Range: 20 uV
@END Instrument  Changes:
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   4.381          6.193          -0.906         Coercive Field: Field at which M//H changes sign
Ms  emu                                 4.155E-4       -4.211E-4      4.183E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -3.471E-6      -3.856E-6      -1.925E-7      Remanent Magnetization: M at H=0        
S                                       0.008          0.009          0.009          Squareness: Mr/Ms                       
S*                                      0.115          0.082          0.098          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
