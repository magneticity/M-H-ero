@Filename: c:\vsm-lv\Will\data\AJA335e-FePtFeRh_1030nm_Tann_6\AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_70deg.VHD
@Measurement Controlfilename: C:\vsm-lv\Will\Recipes\10kOe OoP loop 70deg.VHC
@Signal Manipulation filename: c:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA335e-FePtFeRh_1030nm_Tann_600C
@Date: 05 November 2019    (2019-05-11)
@Time: 15:26:01
@Test ID: AJA335e_FePt_FeRh_Pt_600deg_annealed_OoP_70deg
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 90.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Sample Temperature to 70.0778 [degC] and wait 60.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Applied Field to 9999.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 3:      Set Auto Range Signal to 12.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 5
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 5.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 10000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To: 50.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: 50.0000 [Oe] To: -50.0000 [Oe] Min Stepsize/Sweeprate =  2.0000 [Oe] Max Stepsize/Sweeprate =  2.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -50.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -10000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 4 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 20 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.706
@Y Coils Correction Factor: 0.964
@Sample Shape Correction Factor: 0.919
@Coil Angle Alpha: 42.300
@Coil Angle Beta: -47.320
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
15000.000000   1.000000
15249.000000   1.000524
15499.000000   1.000702
15750.000000   1.001233
16000.000000   1.001406
16250.000000   1.001585
16499.000000   1.001758
16749.000000   1.001937
16999.000000   1.002110
17249.000000   1.001937
17499.000000   1.002289
17749.000000   1.002289
17999.000000   1.002289
18249.000000   1.002462
18499.000000   1.002462
18748.000000   1.002462
18999.000000   1.002462
19249.000000   1.002462
19499.000000   1.002642
19749.000000   1.002642
19999.000000   1.002462
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = No
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 25 October 2019  12:02:56
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 5
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 15:26:01
@@Data
New Section: Section 0: 
2.966600E+1   7.006619E+1   7.006619E+1   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -1.408430E-1   2.347680E-1   -2.399777E-4   -4.931279E-5   4.931279E-5   -2.399777E-4   2.449919E-4   -1.683880E+2   -7.838798E+1   
5.499900E+1   7.002059E+1   7.002059E+1   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -1.239403E-1   2.157549E-1   -2.171445E-4   -4.938433E-5   4.938433E-5   -2.171445E-4   2.226894E-4   -1.671874E+2   -7.718738E+1   
8.010000E+1   7.000399E+1   7.000399E+1   8.998000E+3   8.998000E+3   9.000000E+1   8.998000E+3   8.998000E+3   -1.109894E-1   1.954798E-1   -1.959327E-4   -4.570799E-5   4.570799E-5   -1.959327E-4   2.011936E-4   -1.668687E+2   -7.686865E+1   
1.052490E+2   7.004101E+1   7.004101E+1   8.498000E+3   8.498000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -9.857338E-2   1.780312E-1   -1.768925E-4   -4.348384E-5   4.348384E-5   -1.768925E-4   1.821587E-4   -1.661893E+2   -7.618935E+1   
1.311650E+2   7.004809E+1   7.004809E+1   7.999000E+3   7.999000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -8.703253E-2   1.591426E-1   -1.574555E-4   -3.967098E-5   3.967098E-5   -1.574555E-4   1.623762E-4   -1.658586E+2   -7.585862E+1   
1.569740E+2   7.004699E+1   7.004699E+1   7.498000E+3   7.498000E+3   9.000000E+1   7.498000E+3   7.498000E+3   -7.173275E-2   1.393729E-1   -1.351206E-4   -3.806229E-5   3.806229E-5   -1.351206E-4   1.403792E-4   -1.642679E+2   -7.426794E+1   
1.818330E+2   7.002899E+1   7.002899E+1   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -5.650663E-2   1.205067E-1   -1.134198E-4   -3.698981E-5   3.698981E-5   -1.134198E-4   1.192992E-4   -1.619372E+2   -7.193720E+1   
2.074810E+2   6.998321E+1   6.998321E+1   6.498000E+3   6.498000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -4.784276E-2   1.042727E-1   -9.749035E-5   -3.278458E-5   3.278458E-5   -9.749035E-5   1.028552E-4   -1.614130E+2   -7.141296E+1   
2.323690E+2   6.997979E+1   6.997979E+1   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -3.719939E-2   8.642996E-2   -7.928932E-5   -2.899164E-5   2.899164E-5   -7.928932E-5   8.442340E-5   -1.599154E+2   -6.991538E+1   
2.582520E+2   7.004611E+1   7.004611E+1   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -2.390725E-2   6.874458E-2   -5.955320E-5   -2.726072E-5   2.726072E-5   -5.955320E-5   6.549603E-5   -1.554039E+2   -6.540387E+1   
2.840900E+2   7.002310E+1   7.002310E+1   4.997000E+3   4.997000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -1.104091E-2   5.038763E-2   -3.964294E-5   -2.477581E-5   2.477581E-5   -3.964294E-5   4.674830E-5   -1.479957E+2   -5.799568E+1   
3.096480E+2   7.001119E+1   7.001119E+1   4.498000E+3   4.498000E+3   9.000000E+1   4.498000E+3   4.498000E+3   -2.997377E-4   3.561052E-2   -2.337806E-5   -2.305946E-5   2.305946E-5   -2.337806E-5   3.283706E-5   -1.353931E+2   -4.539310E+1   
3.354910E+2   7.004751E+1   7.004751E+1   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   1.654388E-2   1.447486E-2   8.008780E-7   -2.169962E-5   2.169962E-5   8.008780E-7   2.171440E-5   -8.788632E+1   2.113682E+0   
3.609040E+2   7.002719E+1   7.002719E+1   3.498000E+3   3.498000E+3   9.000000E+1   3.498000E+3   3.498000E+3   2.231468E-2   8.068662E-5   1.374343E-5   -1.655738E-5   1.655738E-5   1.374343E-5   2.151810E-5   -5.030568E+1   3.969432E+1   
3.862030E+2   7.005279E+1   7.005279E+1   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   3.395291E-2   -1.748543E-2   3.237935E-5   -1.368115E-5   1.368115E-5   3.237935E-5   3.515105E-5   -2.290537E+1   6.709463E+1   
4.115470E+2   7.000350E+1   7.000350E+1   2.498000E+3   2.498000E+3   9.000000E+1   2.498000E+3   2.498000E+3   4.796333E-2   -3.413055E-2   5.188204E-5   -1.316158E-5   1.316158E-5   5.188204E-5   5.352544E-5   -1.423466E+1   7.576534E+1   
4.373610E+2   7.001440E+1   7.001440E+1   1.999000E+3   1.999000E+3   9.000000E+1   1.999000E+3   1.999000E+3   5.989149E-2   -5.400444E-2   7.220024E-5   -8.991024E-6   8.991024E-6   7.220024E-5   7.275791E-5   -7.098444E+0   8.290156E+1   
4.714850E+2   7.001980E+1   7.001980E+1   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   6.033234E-2   -5.367524E-2   7.225839E-5   -9.532315E-6   9.532315E-6   7.225839E-5   7.288443E-5   -7.515055E+0   8.248494E+1   
4.937040E+2   7.002770E+1   7.002770E+1   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   6.242067E-2   -5.541724E-2   7.468403E-5   -9.938041E-6   9.938041E-6   7.468403E-5   7.534235E-5   -7.579695E+0   8.242030E+1   
5.160280E+2   6.997949E+1   6.997949E+1   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   6.260628E-2   -5.619402E-2   7.530470E-5   -9.567483E-6   9.567483E-6   7.530470E-5   7.591005E-5   -7.240652E+0   8.275935E+1   
5.382790E+2   7.001339E+1   7.001339E+1   1.799000E+3   1.799000E+3   9.000000E+1   1.799000E+3   1.799000E+3   6.602181E-2   -5.936993E-2   7.948478E-5   -1.001740E-5   1.001740E-5   7.948478E-5   8.011354E-5   -7.183066E+0   8.281693E+1   
5.605560E+2   6.998330E+1   6.998330E+1   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   6.561131E-2   -6.066828E-2   8.007659E-5   -8.864955E-6   8.864955E-6   8.007659E-5   8.056580E-5   -6.317260E+0   8.368274E+1   
5.828390E+2   7.002099E+1   7.002099E+1   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   6.637493E-2   -6.394945E-2   8.268568E-5   -7.284619E-6   7.284619E-6   8.268568E-5   8.300595E-5   -5.034766E+0   8.496523E+1   
6.051230E+2   7.002120E+1   7.002120E+1   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   6.769199E-2   -6.352148E-2   8.322122E-5   -8.538551E-6   8.538551E-6   8.322122E-5   8.365810E-5   -5.858086E+0   8.414191E+1   
6.274070E+2   7.005251E+1   7.005251E+1   1.599000E+3   1.599000E+3   9.000000E+1   1.599000E+3   1.599000E+3   6.931001E-2   -6.552819E-2   8.552851E-5   -8.423351E-6   8.423351E-6   8.552851E-5   8.594230E-5   -5.624687E+0   8.437531E+1   
6.496980E+2   6.998840E+1   6.998840E+1   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   7.042703E-2   -6.859764E-2   8.821820E-5   -7.242815E-6   7.242815E-6   8.821820E-5   8.851502E-5   -4.693522E+0   8.530648E+1   
6.718790E+2   7.000079E+1   7.000079E+1   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   7.195577E-2   -6.796566E-2   8.875174E-5   -8.786693E-6   8.786693E-6   8.875174E-5   8.918563E-5   -5.654032E+0   8.434597E+1   
6.941960E+2   7.002270E+1   7.002270E+1   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   7.092373E-2   -7.112961E-2   9.017433E-5   -5.954864E-6   5.954864E-6   9.017433E-5   9.037074E-5   -3.778169E+0   8.622183E+1   
7.164710E+2   6.999771E+1   6.999771E+1   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   7.436779E-2   -7.221042E-2   9.300753E-5   -7.795592E-6   7.795592E-6   9.300753E-5   9.333366E-5   -4.791149E+0   8.520885E+1   
7.387100E+2   6.998901E+1   6.998901E+1   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   7.414689E-2   -7.448070E-2   9.434956E-5   -6.147968E-6   6.147968E-6   9.434956E-5   9.454966E-5   -3.728213E+0   8.627179E+1   
7.609760E+2   7.001711E+1   7.001711E+1   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   7.496082E-2   -7.697584E-2   9.647784E-5   -5.118723E-6   5.118723E-6   9.647784E-5   9.661353E-5   -3.037034E+0   8.696297E+1   
7.832530E+2   6.996801E+1   6.996801E+1   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   7.739953E-2   -7.688257E-2   9.792481E-5   -6.983439E-6   6.983439E-6   9.792481E-5   9.817351E-5   -4.079103E+0   8.592090E+1   
8.055380E+2   7.002609E+1   7.002609E+1   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   7.788149E-2   -7.915714E-2   9.970419E-5   -5.852872E-6   5.852872E-6   9.970419E-5   9.987583E-5   -3.359543E+0   8.664046E+1   
8.277990E+2   7.001681E+1   7.001681E+1   1.148000E+3   1.148000E+3   9.000000E+1   1.149000E+3   1.149000E+3   7.835058E-2   -8.051715E-2   1.008800E-4   -5.310685E-6   5.310685E-6   1.008800E-4   1.010196E-4   -3.013475E+0   8.698652E+1   
8.500820E+2   7.003280E+1   7.003280E+1   1.098000E+3   1.098000E+3   9.000000E+1   1.099000E+3   1.099000E+3   7.958939E-2   -8.159707E-2   1.023492E-4   -5.520927E-6   5.520927E-6   1.023492E-4   1.024980E-4   -3.087660E+0   8.691234E+1   
8.723340E+2   7.001669E+1   7.001669E+1   1.048000E+3   1.048000E+3   9.000000E+1   1.048000E+3   1.048000E+3   8.107856E-2   -8.478832E-2   1.053483E-4   -4.536011E-6   4.536011E-6   1.053483E-4   1.054459E-4   -2.465477E+0   8.753452E+1   
8.945180E+2   7.003561E+1   7.003561E+1   9.970000E+2   9.970000E+2   9.000000E+1   9.990000E+2   9.990000E+2   8.264536E-2   -8.458830E-2   1.061867E-4   -5.825633E-6   5.825633E-6   1.061867E-4   1.063464E-4   -3.140223E+0   8.685978E+1   
9.163900E+2   7.001171E+1   7.001171E+1   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   8.355715E-2   -8.689535E-2   1.082530E-4   -4.991734E-6   4.991734E-6   1.082530E-4   1.083680E-4   -2.640139E+0   8.735986E+1   
9.382410E+2   7.001821E+1   7.001821E+1   8.980000E+2   8.980000E+2   9.000000E+1   8.990000E+2   8.990000E+2   8.365870E-2   -8.766818E-2   1.088191E-4   -4.561598E-6   4.561598E-6   1.088191E-4   1.089146E-4   -2.400382E+0   8.759962E+1   
9.601660E+2   7.003631E+1   7.003631E+1   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   8.528010E-2   -9.081681E-2   1.118722E-4   -3.702347E-6   3.702347E-6   1.118722E-4   1.119334E-4   -1.895480E+0   8.810452E+1   
9.819850E+2   7.002181E+1   7.002181E+1   7.980000E+2   7.980000E+2   9.000000E+1   7.980000E+2   7.980000E+2   8.635694E-2   -9.049898E-2   1.123309E-4   -4.706605E-6   4.706605E-6   1.123309E-4   1.124295E-4   -2.399259E+0   8.760074E+1   
1.003848E+3   7.007031E+1   7.007031E+1   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   8.742335E-2   -9.356948E-2   1.149900E-4   -3.487946E-6   3.487946E-6   1.149900E-4   1.150429E-4   -1.737397E+0   8.826260E+1   
1.025667E+3   7.000350E+1   7.000350E+1   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   8.809276E-2   -9.479241E-2   1.162004E-4   -3.183542E-6   3.183542E-6   1.162004E-4   1.162440E-4   -1.569341E+0   8.843066E+1   
1.047544E+3   7.002279E+1   7.002279E+1   6.480000E+2   6.480000E+2   9.000000E+1   6.480000E+2   6.480000E+2   8.880454E-2   -9.581195E-2   1.173044E-4   -3.043450E-6   3.043450E-6   1.173044E-4   1.173439E-4   -1.486199E+0   8.851380E+1   
1.069364E+3   7.004559E+1   7.004559E+1   5.980000E+2   5.980000E+2   9.000000E+1   5.990000E+2   5.990000E+2   9.022377E-2   -9.738768E-2   1.192081E-4   -3.062985E-6   3.062985E-6   1.192081E-4   1.192475E-4   -1.471859E+0   8.852814E+1   
1.091240E+3   7.004629E+1   7.004629E+1   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   9.294694E-2   -9.913552E-2   1.220301E-4   -3.934440E-6   3.934440E-6   1.220301E-4   1.220935E-4   -1.846666E+0   8.815333E+1   
1.113126E+3   7.002499E+1   7.002499E+1   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   9.290983E-2   -1.002857E-1   1.227562E-4   -3.155045E-6   3.155045E-6   1.227562E-4   1.227968E-4   -1.472275E+0   8.852772E+1   
1.135006E+3   7.004571E+1   7.004571E+1   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   9.241741E-2   -1.032383E-1   1.243748E-4   -8.605217E-7   8.605217E-7   1.243748E-4   1.243777E-4   -3.964106E-1   8.960359E+1   
1.156880E+3   7.000839E+1   7.000839E+1   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   9.428341E-2   -1.039418E-1   1.259866E-4   -1.780760E-6   1.780760E-6   1.259866E-4   1.259992E-4   -8.097945E-1   8.919021E+1   
1.178706E+3   7.001910E+1   7.001910E+1   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   9.615065E-2   -1.053091E-1   1.280315E-4   -2.267882E-6   2.267882E-6   1.280315E-4   1.280516E-4   -1.014801E+0   8.898520E+1   
1.200530E+3   7.005020E+1   7.005020E+1   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   9.779419E-2   -1.058595E-1   1.294061E-4   -3.123664E-6   3.123664E-6   1.294061E-4   1.294438E-4   -1.382763E+0   8.861724E+1   
1.222412E+3   7.001959E+1   7.001959E+1   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   9.653049E-2   -1.078954E-1   1.299508E-4   -8.580070E-7   8.580070E-7   1.299508E-4   1.299536E-4   -3.782930E-1   8.962171E+1   
1.244293E+3   7.001199E+1   7.001199E+1   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   9.796905E-2   -1.091532E-1   1.316594E-4   -1.099669E-6   1.099669E-6   1.316594E-4   1.316640E-4   -4.785450E-1   8.952146E+1   
1.266173E+3   7.004290E+1   7.004290E+1   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   9.912876E-2   -1.122261E-1   1.343777E-4   5.151100E-8   -5.151100E-8   1.343777E-4   1.343777E-4   2.196319E-2   9.002196E+1   
1.287979E+3   7.001730E+1   7.001730E+1   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   1.006305E-1   -1.124531E-1   1.354540E-4   -9.108052E-7   9.108052E-7   1.354540E-4   1.354571E-4   -3.852563E-1   8.961474E+1   
1.309667E+3   7.005261E+1   7.005261E+1   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   1.017285E-1   -1.136720E-1   1.369267E-4   -9.260459E-7   9.260459E-7   1.369267E-4   1.369298E-4   -3.874899E-1   8.961251E+1   
1.342838E+3   7.005660E+1   7.005660E+1   4.700000E+1   4.700000E+1   9.000000E+1   4.700000E+1   4.700000E+1   1.012269E-1   -1.150126E-1   1.374897E-4   3.214403E-7   -3.214403E-7   1.374897E-4   1.374901E-4   1.339528E-1   9.013395E+1   
1.364188E+3   7.000680E+1   7.000680E+1   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   1.014411E-1   -1.141631E-1   1.370688E-4   -3.923232E-7   3.923232E-7   1.370688E-4   1.370694E-4   -1.639935E-1   8.983601E+1   
1.383197E+3   6.998910E+1   6.998910E+1   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   1.017828E-1   -1.143705E-1   1.374152E-4   -5.095227E-7   5.095227E-7   1.374152E-4   1.374162E-4   -2.124464E-1   8.978755E+1   
1.405605E+3   7.000451E+1   7.000451E+1   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   1.033475E-1   -1.135045E-1   1.378185E-4   -2.232983E-6   2.232983E-6   1.378185E-4   1.378366E-4   -9.282451E-1   8.907175E+1   
1.424682E+3   7.002160E+1   7.002160E+1   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   1.027394E-1   -1.142674E-1   1.379395E-4   -1.284426E-6   1.284426E-6   1.379395E-4   1.379455E-4   -5.334955E-1   8.946650E+1   
1.447108E+3   7.003671E+1   7.003671E+1   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   1.016724E-1   -1.145555E-1   1.374674E-4   -3.068906E-7   3.068906E-7   1.374674E-4   1.374678E-4   -1.279104E-1   8.987209E+1   
1.466242E+3   7.002200E+1   7.002200E+1   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   1.015727E-1   -1.150114E-1   1.377027E-4   6.491344E-8   -6.491344E-8   1.377027E-4   1.377027E-4   2.700939E-2   9.002701E+1   
1.488669E+3   6.997970E+1   6.997970E+1   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   1.007014E-1   -1.146706E-1   1.369420E-4   4.865028E-7   -4.865028E-7   1.369420E-4   1.369429E-4   2.035492E-1   9.020355E+1   
1.507789E+3   7.001010E+1   7.001010E+1   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   1.022363E-1   -1.142484E-1   1.376160E-4   -9.247178E-7   9.247178E-7   1.376160E-4   1.376191E-4   -3.849960E-1   8.961500E+1   
1.530222E+3   7.004180E+1   7.004180E+1   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   1.016193E-1   -1.135382E-1   1.367720E-4   -9.327389E-7   9.327389E-7   1.367720E-4   1.367752E-4   -3.907318E-1   8.960927E+1   
1.549287E+3   6.995730E+1   6.995730E+1   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   1.029943E-1   -1.143543E-1   1.381536E-4   -1.416211E-6   1.416211E-6   1.381536E-4   1.381609E-4   -5.873174E-1   8.941268E+1   
1.571683E+3   7.002621E+1   7.002621E+1   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   1.025765E-1   -1.144423E-1   1.379527E-4   -1.049612E-6   1.049612E-6   1.379527E-4   1.379567E-4   -4.359261E-1   8.956407E+1   
1.590656E+3   7.000649E+1   7.000649E+1   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   1.015309E-1   -1.151461E-1   1.377646E-4   1.838221E-7   -1.838221E-7   1.377646E-4   1.377647E-4   7.645086E-2   9.007645E+1   
1.612992E+3   7.001019E+1   7.001019E+1   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   1.036463E-1   -1.136913E-1   1.381249E-4   -2.331857E-6   2.331857E-6   1.381249E-4   1.381446E-4   -9.671888E-1   8.903281E+1   
1.632064E+3   7.001821E+1   7.001821E+1   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   1.020816E-1   -1.146933E-1   1.378102E-4   -5.195077E-7   5.195077E-7   1.378102E-4   1.378111E-4   -2.159888E-1   8.978401E+1   
1.654489E+3   6.998571E+1   6.998571E+1   1.700000E+1   1.700000E+1   9.000000E+1   1.700000E+1   1.700000E+1   1.011152E-1   -1.164073E-1   1.383290E-4   1.315841E-6   -1.315841E-6   1.383290E-4   1.383353E-4   5.450039E-1   9.054500E+1   
1.675834E+3   6.998611E+1   6.998611E+1   1.500000E+1   1.500000E+1   9.000000E+1   1.500000E+1   1.500000E+1   1.027106E-1   -1.139926E-1   1.377426E-4   -1.442810E-6   1.442810E-6   1.377426E-4   1.377502E-4   -6.001329E-1   8.939987E+1   
1.697210E+3   7.005251E+1   7.005251E+1   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   1.036288E-1   -1.150034E-1   1.389687E-4   -1.461083E-6   1.461083E-6   1.389687E-4   1.389764E-4   -6.023719E-1   8.939763E+1   
1.716220E+3   7.003591E+1   7.003591E+1   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   1.025943E-1   -1.151004E-1   1.383923E-4   -6.325452E-7   6.325452E-7   1.383923E-4   1.383937E-4   -2.618782E-1   8.973812E+1   
1.738301E+3   7.004669E+1   7.004669E+1   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   1.014524E-1   -1.152268E-1   1.377686E-4   2.946583E-7   -2.946583E-7   1.377686E-4   1.377689E-4   1.225435E-1   9.012254E+1   
1.757041E+3   7.003100E+1   7.003100E+1   9.000000E+0   9.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   1.024924E-1   -1.150528E-1   1.382983E-4   -5.882920E-7   5.882920E-7   1.382983E-4   1.382996E-4   -2.437228E-1   8.975628E+1   
1.778723E+3   7.003890E+1   7.003890E+1   5.000000E+0   5.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   1.026219E-1   -1.157459E-1   1.388297E-4   -2.309489E-7   2.309489E-7   1.388297E-4   1.388299E-4   -9.531379E-2   8.990469E+1   
1.799809E+3   7.002700E+1   7.002700E+1   3.000000E+0   3.000000E+0   9.000000E+1   3.000000E+0   3.000000E+0   1.036908E-1   -1.146647E-1   1.387864E-4   -1.728344E-6   1.728344E-6   1.387864E-4   1.387972E-4   -7.134827E-1   8.928652E+1   
1.820840E+3   7.003951E+1   7.003951E+1   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   1.025397E-1   -1.157229E-1   1.387639E-4   -1.851958E-7   1.851958E-7   1.387639E-4   1.387640E-4   -7.646751E-2   8.992353E+1   
1.839520E+3   7.001550E+1   7.001550E+1   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   1.016653E-1   -1.162659E-1   1.385770E-4   8.165271E-7   -8.165271E-7   1.385770E-4   1.385794E-4   3.375958E-1   9.033760E+1   
1.861500E+3   7.000680E+1   7.000680E+1   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   1.020482E-1   -1.160183E-1   1.386525E-4   3.714819E-7   -3.714819E-7   1.386525E-4   1.386530E-4   1.535082E-1   9.015351E+1   
1.883543E+3   7.003329E+1   7.003329E+1   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   1.030253E-1   -1.152354E-1   1.387467E-4   -8.631045E-7   8.631045E-7   1.387467E-4   1.387493E-4   -3.564165E-1   8.964358E+1   
1.905551E+3   7.003631E+1   7.003631E+1   -5.000000E+0   -5.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   1.031235E-1   -1.156624E-1   1.390855E-4   -6.565249E-7   6.565249E-7   1.390855E-4   1.390871E-4   -2.704511E-1   8.972955E+1   
1.927319E+3   7.000970E+1   7.000970E+1   -8.000000E+0   -8.000000E+0   9.000000E+1   -6.000000E+0   -6.000000E+0   1.045286E-1   -1.148332E-1   1.394141E-4   -2.237925E-6   2.237925E-6   1.394141E-4   1.394321E-4   -9.196532E-1   8.908035E+1   
1.949506E+3   7.002010E+1   7.002010E+1   -1.000000E+1   -1.000000E+1   9.000000E+1   -8.000000E+0   -8.000000E+0   1.026624E-1   -1.152679E-1   1.385435E-4   -5.734001E-7   5.734001E-7   1.385435E-4   1.385447E-4   -2.371329E-1   8.976287E+1   
1.971651E+3   7.005319E+1   7.005319E+1   -1.100000E+1   -1.100000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   1.026241E-1   -1.162088E-1   1.391326E-4   7.012104E-8   -7.012104E-8   1.391326E-4   1.391326E-4   2.887634E-2   9.002888E+1   
1.993591E+3   7.005041E+1   7.005041E+1   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   1.033803E-1   -1.156425E-1   1.392313E-4   -8.594937E-7   8.594937E-7   1.392313E-4   1.392339E-4   -3.536902E-1   8.964631E+1   
2.015774E+3   7.001061E+1   7.001061E+1   -1.500000E+1   -1.500000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   1.030800E-1   -1.163791E-1   1.395253E-4   -1.557740E-7   1.557740E-7   1.395253E-4   1.395254E-4   -6.396825E-2   8.993603E+1   
2.037692E+3   7.004901E+1   7.004901E+1   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   1.030333E-1   -1.161352E-1   1.393376E-4   -2.807084E-7   2.807084E-7   1.393376E-4   1.393379E-4   -1.154274E-1   8.988457E+1   
2.059857E+3   7.002450E+1   7.002450E+1   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   1.032732E-1   -1.176029E-1   1.404418E-4   5.013788E-7   -5.013788E-7   1.404418E-4   1.404427E-4   2.045456E-1   9.020455E+1   
2.082101E+3   6.998040E+1   6.998040E+1   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   1.020654E-1   -1.158042E-1   1.385236E-4   2.187662E-7   -2.187662E-7   1.385236E-4   1.385238E-4   9.048542E-2   9.009049E+1   
2.104341E+3   6.999621E+1   6.999621E+1   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   1.026167E-1   -1.162248E-1   1.391384E-4   8.601418E-8   -8.601418E-8   1.391384E-4   1.391384E-4   3.541976E-2   9.003542E+1   
2.126584E+3   7.002361E+1   7.002361E+1   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   1.030238E-1   -1.165813E-1   1.396223E-4   1.794767E-8   -1.794767E-8   1.396223E-4   1.396223E-4   7.365053E-3   9.000737E+1   
2.148823E+3   7.002130E+1   7.002130E+1   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   1.034002E-1   -1.168062E-1   1.400015E-4   -1.134525E-7   1.134525E-7   1.400015E-4   1.400015E-4   -4.643057E-2   8.995357E+1   
2.170996E+3   7.003390E+1   7.003390E+1   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   1.025201E-1   -1.164000E-1   1.391928E-4   2.719894E-7   -2.719894E-7   1.391928E-4   1.391930E-4   1.119586E-1   9.011196E+1   
2.193229E+3   7.003161E+1   7.003161E+1   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   1.033281E-1   -1.164524E-1   1.397265E-4   -2.914023E-7   2.914023E-7   1.397265E-4   1.397268E-4   -1.194912E-1   8.988051E+1   
2.215453E+3   7.005639E+1   7.005639E+1   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   1.034843E-1   -1.174685E-1   1.404849E-4   2.573891E-7   -2.573891E-7   1.404849E-4   1.404851E-4   1.049742E-1   9.010497E+1   
2.237744E+3   7.004730E+1   7.004730E+1   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   1.024673E-1   -1.173081E-1   1.397516E-4   9.047232E-7   -9.047232E-7   1.397516E-4   1.397545E-4   3.709160E-1   9.037092E+1   
2.260009E+3   7.003210E+1   7.003210E+1   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   1.051539E-1   -1.156609E-1   1.403398E-4   -2.159235E-6   2.159235E-6   1.403398E-4   1.403564E-4   -8.814700E-1   8.911853E+1   
2.282272E+3   7.003069E+1   7.003069E+1   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   1.026633E-1   -1.167835E-1   1.395311E-4   4.167451E-7   -4.167451E-7   1.395311E-4   1.395317E-4   1.711279E-1   9.017113E+1   
2.304534E+3   7.002319E+1   7.002319E+1   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   1.034328E-1   -1.186850E-1   1.412452E-4   1.090802E-6   -1.090802E-6   1.412452E-4   1.412494E-4   4.424724E-1   9.044247E+1   
2.326754E+3   7.004711E+1   7.004711E+1   -4.300000E+1   -4.300000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   1.025093E-1   -1.170280E-1   1.395951E-4   6.905025E-7   -6.905025E-7   1.395951E-4   1.395968E-4   2.834093E-1   9.028341E+1   
2.348730E+3   6.999560E+1   6.999560E+1   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   1.028281E-1   -1.172440E-1   1.399329E-4   5.959549E-7   -5.959549E-7   1.399329E-4   1.399341E-4   2.440134E-1   9.024401E+1   
2.371042E+3   7.004189E+1   7.004189E+1   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.600000E+1   -4.600000E+1   1.043648E-1   -1.163297E-1   1.402875E-4   -1.138351E-6   1.138351E-6   1.402875E-4   1.402921E-4   -4.649117E-1   8.953509E+1   
2.393269E+3   7.001751E+1   7.001751E+1   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   1.031594E-1   -1.169022E-1   1.399151E-4   1.274458E-7   -1.274458E-7   1.399151E-4   1.399152E-4   5.218955E-2   9.005219E+1   
2.426609E+3   7.002319E+1   7.002319E+1   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   1.060429E-1   -1.184567E-1   1.427103E-4   -9.890114E-7   9.890114E-7   1.427103E-4   1.427137E-4   -3.970651E-1   8.960293E+1   
2.448284E+3   7.008340E+1   7.008340E+1   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   1.056886E-1   -1.203788E-1   1.437430E-4   5.296758E-7   -5.296758E-7   1.437430E-4   1.437440E-4   2.111271E-1   9.021113E+1   
2.469965E+3   7.000771E+1   7.000771E+1   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   1.065841E-1   -1.218931E-1   1.452830E-4   8.573135E-7   -8.573135E-7   1.452830E-4   1.452855E-4   3.380979E-1   9.033810E+1   
2.491703E+3   7.002691E+1   7.002691E+1   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   1.075478E-1   -1.241514E-1   1.473495E-4   1.620984E-6   -1.620984E-6   1.473495E-4   1.473584E-4   6.302822E-1   9.063028E+1   
2.513895E+3   7.001000E+1   7.001000E+1   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   1.082433E-1   -1.242278E-1   1.478293E-4   1.156536E-6   -1.156536E-6   1.478293E-4   1.478338E-4   4.482417E-1   9.044824E+1   
2.535585E+3   6.998861E+1   6.998861E+1   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   1.096634E-1   -1.251899E-1   1.493339E-4   7.351374E-7   -7.351374E-7   1.493339E-4   1.493357E-4   2.820521E-1   9.028205E+1   
2.557325E+3   7.002429E+1   7.002429E+1   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   1.102331E-1   -1.262109E-1   1.503511E-4   9.812753E-7   -9.812753E-7   1.503511E-4   1.503543E-4   3.739390E-1   9.037394E+1   
2.579512E+3   7.000280E+1   7.000280E+1   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   1.103730E-1   -1.289637E-1   1.522305E-4   2.677548E-6   -2.677548E-6   1.522305E-4   1.522540E-4   1.007659E+0   9.100766E+1   
2.601155E+3   6.999691E+1   6.999691E+1   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   1.128446E-1   -1.306161E-1   1.548347E-4   1.929774E-6   -1.929774E-6   1.548347E-4   1.548467E-4   7.140662E-1   9.071407E+1   
2.622829E+3   7.002410E+1   7.002410E+1   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   1.120018E-1   -1.311407E-1   1.546553E-4   2.896104E-6   -2.896104E-6   1.546553E-4   1.546824E-4   1.072806E+0   9.107281E+1   
2.644516E+3   7.000701E+1   7.000701E+1   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   1.145463E-1   -1.316043E-1   1.565304E-4   1.317157E-6   -1.317157E-6   1.565304E-4   1.565359E-4   4.821156E-1   9.048212E+1   
2.666205E+3   7.005001E+1   7.005001E+1   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.490000E+2   -6.490000E+2   1.138438E-1   -1.347382E-1   1.581371E-4   3.885624E-6   -3.885624E-6   1.581371E-4   1.581848E-4   1.407545E+0   9.140755E+1   
2.687885E+3   7.004791E+1   7.004791E+1   -7.000000E+2   -7.000000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   1.158833E-1   -1.362663E-1   1.603933E-4   3.376173E-6   -3.376173E-6   1.603933E-4   1.604288E-4   1.205860E+0   9.120586E+1   
2.709508E+3   7.000411E+1   7.000411E+1   -7.500000E+2   -7.500000E+2   9.000000E+1   -7.490000E+2   -7.490000E+2   1.165552E-1   -1.367943E-1   1.611526E-4   3.224402E-6   -3.224402E-6   1.611526E-4   1.611848E-4   1.146243E+0   9.114624E+1   
2.731242E+3   7.003149E+1   7.003149E+1   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   1.179891E-1   -1.387338E-1   1.633023E-4   3.431823E-6   -3.431823E-6   1.633023E-4   1.633383E-4   1.203902E+0   9.120390E+1   
2.752956E+3   7.002331E+1   7.002331E+1   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   1.181751E-1   -1.399230E-1   1.641917E-4   4.071741E-6   -4.071741E-6   1.641917E-4   1.642422E-4   1.420570E+0   9.142057E+1   
2.774633E+3   7.000659E+1   7.000659E+1   -9.000000E+2   -9.000000E+2   9.000000E+1   -8.990000E+2   -8.990000E+2   1.195943E-1   -1.418898E-1   1.663501E-4   4.307916E-6   -4.307916E-6   1.663501E-4   1.664059E-4   1.483439E+0   9.148344E+1   
2.796264E+3   7.002941E+1   7.002941E+1   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   1.201161E-1   -1.424344E-1   1.670274E-4   4.277949E-6   -4.277949E-6   1.670274E-4   1.670822E-4   1.467153E+0   9.146715E+1   
2.817972E+3   7.000610E+1   7.000610E+1   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   1.204828E-1   -1.440235E-1   1.682891E-4   5.045739E-6   -5.045739E-6   1.682891E-4   1.683647E-4   1.717360E+0   9.171736E+1   
2.840460E+3   6.998760E+1   6.998760E+1   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   1.222272E-1   -1.453765E-1   1.702488E-4   4.640034E-6   -4.640034E-6   1.702488E-4   1.703120E-4   1.561178E+0   9.156118E+1   
2.862254E+3   7.001660E+1   7.001660E+1   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   1.221624E-1   -1.475443E-1   1.716206E-4   6.105172E-6   -6.105172E-6   1.716206E-4   1.717291E-4   2.037361E+0   9.203736E+1   
2.884122E+3   7.007031E+1   7.007031E+1   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   1.224355E-1   -1.491050E-1   1.728058E-4   6.923514E-6   -6.923514E-6   1.728058E-4   1.729445E-4   2.294344E+0   9.229434E+1   
2.906725E+3   7.000790E+1   7.000790E+1   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   1.236673E-1   -1.500250E-1   1.741666E-4   6.613981E-6   -6.613981E-6   1.741666E-4   1.742921E-4   2.174764E+0   9.217476E+1   
2.928844E+3   7.001199E+1   7.001199E+1   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   1.267588E-1   -1.511675E-1   1.768220E-4   5.074317E-6   -5.074317E-6   1.768220E-4   1.768948E-4   1.643784E+0   9.164378E+1   
2.950734E+3   7.003771E+1   7.003771E+1   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   1.270441E-1   -1.516685E-1   1.773247E-4   5.190815E-6   -5.190815E-6   1.773247E-4   1.774007E-4   1.676737E+0   9.167674E+1   
2.973054E+3   7.002801E+1   7.002801E+1   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   1.273555E-1   -1.544628E-1   1.793371E-4   6.787303E-6   -6.787303E-6   1.793371E-4   1.794655E-4   2.167417E+0   9.216742E+1   
2.995134E+3   7.000430E+1   7.000430E+1   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   1.268297E-1   -1.554593E-1   1.796610E-4   7.827700E-6   -7.827700E-6   1.796610E-4   1.798314E-4   2.494758E+0   9.249476E+1   
3.017252E+3   7.005349E+1   7.005349E+1   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   1.299402E-1   -1.571816E-1   1.827058E-4   6.653038E-6   -6.653038E-6   1.827058E-4   1.828269E-4   2.085443E+0   9.208544E+1   
3.039594E+3   7.001940E+1   7.001940E+1   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   1.295954E-1   -1.589892E-1   1.836699E-4   8.089861E-6   -8.089861E-6   1.836699E-4   1.838480E-4   2.522000E+0   9.252200E+1   
3.061614E+3   7.000421E+1   7.000421E+1   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.548000E+3   -1.548000E+3   1.305861E-1   -1.591472E-1   1.843853E-4   7.460451E-6   -7.460451E-6   1.843853E-4   1.845362E-4   2.316992E+0   9.231699E+1   
3.084192E+3   7.002050E+1   7.002050E+1   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   1.319915E-1   -1.612813E-1   1.866441E-4   7.816151E-6   -7.816151E-6   1.866441E-4   1.868077E-4   2.397992E+0   9.239799E+1   
3.107040E+3   7.000390E+1   7.000390E+1   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   1.349907E-1   -1.634153E-1   1.898882E-4   6.993021E-6   -6.993021E-6   1.898882E-4   1.900169E-4   2.109081E+0   9.210908E+1   
3.128847E+3   6.999151E+1   6.999151E+1   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.698000E+3   -1.698000E+3   1.341261E-1   -1.632199E-1   1.892264E-4   7.504707E-6   -7.504707E-6   1.892264E-4   1.893752E-4   2.271156E+0   9.227116E+1   
3.150952E+3   7.001281E+1   7.001281E+1   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.748000E+3   -1.748000E+3   1.339319E-1   -1.661099E-1   1.909886E-4   9.537728E-6   -9.537728E-6   1.909886E-4   1.912266E-4   2.858904E+0   9.285890E+1   
3.174586E+3   7.000320E+1   7.000320E+1   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.798000E+3   -1.798000E+3   1.354769E-1   -1.669606E-1   1.924978E-4   8.951169E-6   -8.951169E-6   1.924978E-4   1.927058E-4   2.662342E+0   9.266234E+1   
3.197154E+3   7.002691E+1   7.002691E+1   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.848000E+3   -1.848000E+3   1.368532E-1   -1.689588E-1   1.946501E-4   9.239570E-6   -9.239570E-6   1.946501E-4   1.948693E-4   2.717652E+0   9.271765E+1   
3.219465E+3   6.999471E+1   6.999471E+1   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   1.366851E-1   -1.696730E-1   1.950113E-4   9.830855E-6   -9.830855E-6   1.950113E-4   1.952590E-4   2.885935E+0   9.288594E+1   
3.242809E+3   7.000302E+1   7.000302E+1   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   1.391094E-1   -1.723037E-1   1.982235E-4   9.757672E-6   -9.757672E-6   1.982235E-4   1.984635E-4   2.818145E+0   9.281814E+1   
3.265098E+3   6.998730E+1   6.998730E+1   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   1.387415E-1   -1.723065E-1   1.979979E-4   1.003154E-5   -1.003154E-5   1.979979E-4   1.982518E-4   2.900406E+0   9.290041E+1   
3.302090E+3   7.003631E+1   7.003631E+1   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.466850E-1   -1.887027E-1   2.135876E-4   1.487572E-5   -1.487572E-5   2.135876E-4   2.141050E-4   3.984042E+0   9.398404E+1   
3.328282E+3   7.002590E+1   7.002590E+1   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.575194E-1   -2.031561E-1   2.296993E-4   1.631149E-5   -1.631149E-5   2.296993E-4   2.302777E-4   4.061890E+0   9.406189E+1   
3.353442E+3   6.999481E+1   6.999481E+1   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.675481E-1   -2.195112E-1   2.465514E-4   1.958642E-5   -1.958642E-5   2.465514E-4   2.473282E-4   4.542125E+0   9.454212E+1   
3.379091E+3   7.003188E+1   7.003188E+1   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   1.753106E-1   -2.346815E-1   2.612307E-4   2.376299E-5   -2.376299E-5   2.612307E-4   2.623093E-4   5.197635E+0   9.519763E+1   
3.404878E+3   7.001629E+1   7.001629E+1   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   1.825997E-1   -2.476661E-1   2.741940E-4   2.686072E-5   -2.686072E-5   2.741940E-4   2.755065E-4   5.594985E+0   9.559498E+1   
3.429607E+3   7.001650E+1   7.001650E+1   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   1.866732E-1   -2.561481E-1   2.822366E-4   2.939309E-5   -2.939309E-5   2.822366E-4   2.837630E-4   5.945547E+0   9.594555E+1   
3.454846E+3   6.998919E+1   6.998919E+1   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   1.854729E-1   -2.568195E-1   2.819318E-4   3.071986E-5   -3.071986E-5   2.819318E-4   2.836006E-4   6.218531E+0   9.621853E+1   
3.481043E+3   7.003491E+1   7.003491E+1   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   1.722120E-1   -2.442816E-1   2.655675E-4   3.233112E-5   -3.233112E-5   2.655675E-4   2.675283E-4   6.941230E+0   9.694123E+1   
3.506191E+3   7.004601E+1   7.004601E+1   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.503751E-1   -2.233449E-1   2.384311E-4   3.479449E-5   -3.479449E-5   2.384311E-4   2.409565E-4   8.302626E+0   9.830263E+1   
3.530889E+3   7.002130E+1   7.002130E+1   -7.000000E+3   -7.000000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.298093E-1   -2.026597E-1   2.122443E-4   3.648224E-5   -3.648224E-5   2.122443E-4   2.153569E-4   9.753147E+0   9.975315E+1   
3.556091E+3   6.997811E+1   6.997811E+1   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.177504E-1   -1.913834E-1   1.974448E-4   3.802920E-5   -3.802920E-5   1.974448E-4   2.010738E-4   1.090205E+1   1.009020E+2   
3.581285E+3   7.002371E+1   7.002371E+1   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.129814E-1   -1.892167E-1   1.930852E-4   4.013999E-5   -4.013999E-5   1.930852E-4   1.972134E-4   1.174380E+1   1.017438E+2   
3.606947E+3   7.004089E+1   7.004089E+1   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.116778E-1   -1.907394E-1   1.932710E-4   4.209963E-5   -4.209963E-5   1.932710E-4   1.978030E-4   1.228861E+1   1.022886E+2   
3.632663E+3   7.001180E+1   7.001180E+1   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.098453E-1   -1.952939E-1   1.951044E-4   4.643260E-5   -4.643260E-5   1.951044E-4   2.005535E-4   1.338671E+1   1.033867E+2   
3.658346E+3   7.004940E+1   7.004940E+1   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.202784E-1   -2.106590E-1   2.115617E-4   4.876125E-5   -4.876125E-5   2.115617E-4   2.171083E-4   1.297901E+1   1.029790E+2   
3.683587E+3   7.004711E+1   7.004711E+1   -9.999000E+3   -9.999000E+3   9.000000E+1   -9.998000E+3   -9.998000E+3   1.280974E-1   -2.227506E-1   2.242709E-4   5.088329E-5   -5.088329E-5   2.242709E-4   2.299707E-4   1.278304E+1   1.027830E+2   
3.720161E+3   7.003329E+1   7.003329E+1   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.164754E-1   -2.039795E-1   2.048602E-4   4.720721E-5   -4.720721E-5   2.048602E-4   2.102290E-4   1.297650E+1   1.029765E+2   
3.744352E+3   7.002599E+1   7.002599E+1   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.031514E-1   -1.881364E-1   1.863042E-4   4.670428E-5   -4.670428E-5   1.863042E-4   1.920691E-4   1.407335E+1   1.040734E+2   
3.768589E+3   7.002090E+1   7.002090E+1   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   9.299543E-2   -1.713508E-1   1.690931E-4   4.324202E-5   -4.324202E-5   1.690931E-4   1.745347E-4   1.434477E+1   1.043448E+2   
3.793194E+3   7.001681E+1   7.001681E+1   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   8.542459E-2   -1.549981E-1   1.537621E-4   3.815072E-5   -3.815072E-5   1.537621E-4   1.584243E-4   1.393456E+1   1.039346E+2   
3.817890E+3   7.002001E+1   7.002001E+1   -7.499000E+3   -7.499000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   7.302772E-2   -1.395321E-1   1.360249E-4   3.720858E-5   -3.720858E-5   1.360249E-4   1.410222E-4   1.529858E+1   1.052986E+2   
3.843082E+3   7.002120E+1   7.002120E+1   -7.000000E+3   -7.000000E+3   9.000000E+1   -6.999000E+3   -6.999000E+3   6.384942E-2   -1.242465E-1   1.203951E-4   3.400384E-5   -3.400384E-5   1.203951E-4   1.251049E-4   1.577155E+1   1.057716E+2   
3.867818E+3   6.998010E+1   6.998010E+1   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   5.525860E-2   -1.083629E-1   1.047391E-4   2.997364E-5   -2.997364E-5   1.047391E-4   1.089435E-4   1.596977E+1   1.059698E+2   
3.891968E+3   6.998910E+1   6.998910E+1   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   4.572522E-2   -9.441532E-2   8.976117E-5   2.790628E-5   -2.790628E-5   8.976117E-5   9.399909E-5   1.727019E+1   1.072702E+2   
3.916641E+3   7.002191E+1   7.002191E+1   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   3.577283E-2   -7.742805E-2   7.254450E-5   2.416158E-5   -2.416158E-5   7.254450E-5   7.646232E-5   1.842079E+1   1.084208E+2   
3.941778E+3   7.001959E+1   7.001959E+1   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   2.380816E-2   -5.952179E-2   5.348523E-5   2.130441E-5   -2.130441E-5   5.348523E-5   5.757211E-5   2.171854E+1   1.117185E+2   
3.966531E+3   7.001089E+1   7.001089E+1   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   1.412972E-2   -4.569976E-2   3.849942E-5   1.942643E-5   -1.942643E-5   3.849942E-5   4.312298E-5   2.677507E+1   1.167751E+2   
3.991165E+3   7.002819E+1   7.002819E+1   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   6.938458E-3   -2.984620E-2   2.372819E-5   1.438070E-5   -1.438070E-5   2.372819E-5   2.774584E-5   3.121837E+1   1.212184E+2   
4.015841E+3   7.005670E+1   7.005670E+1   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   -6.374264E-3   -1.359835E-2   4.915593E-6   1.360482E-5   -1.360482E-5   4.915593E-6   1.446562E-5   7.013458E+1   1.601346E+2   
4.040030E+3   7.001809E+1   7.001809E+1   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   -1.485651E-2   7.998124E-4   -9.705899E-6   1.046544E-5   -1.046544E-5   -9.705899E-6   1.427340E-5   1.328436E+2   2.228436E+2   
4.064766E+3   7.002529E+1   7.002529E+1   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   -2.441623E-2   1.874635E-2   -2.730455E-5   5.803170E-6   -5.803170E-6   -2.730455E-5   2.791443E-5   1.680012E+2   2.580012E+2   
4.089420E+3   7.005181E+1   7.005181E+1   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   -3.460117E-2   3.368479E-2   -4.333061E-5   3.569940E-6   -3.569940E-6   -4.333061E-5   4.347742E-5   1.752901E+2   2.652901E+2   
4.123082E+3   7.000302E+1   7.000302E+1   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.948000E+3   -1.948000E+3   -3.453152E-2   3.762859E-2   -4.585610E-5   9.400709E-7   -9.400709E-7   -4.585610E-5   4.586574E-5   1.788256E+2   2.688256E+2   
4.144857E+3   7.004669E+1   7.004669E+1   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   -3.637413E-2   3.899322E-2   -4.788406E-5   1.410772E-6   -1.410772E-6   -4.788406E-5   4.790483E-5   1.783124E+2   2.683124E+2   
4.166956E+3   6.999819E+1   6.999819E+1   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.849000E+3   -1.849000E+3   -3.733193E-2   4.010534E-2   -4.920053E-5   1.392120E-6   -1.392120E-6   -4.920053E-5   4.922022E-5   1.783793E+2   2.683793E+2   
4.188799E+3   7.006039E+1   7.006039E+1   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.798000E+3   -1.798000E+3   -3.874625E-2   4.193873E-2   -5.126900E-5   1.239572E-6   -1.239572E-6   -5.126900E-5   5.128398E-5   1.786150E+2   2.686150E+2   
4.210592E+3   7.003079E+1   7.003079E+1   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   -3.970989E-2   4.230563E-2   -5.210372E-5   1.712439E-6   -1.712439E-6   -5.210372E-5   5.213185E-5   1.781176E+2   2.681176E+2   
4.232684E+3   6.996191E+1   6.996191E+1   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   -4.134202E-2   4.456520E-2   -5.458441E-5   1.442380E-6   -1.442380E-6   -5.458441E-5   5.460347E-5   1.784863E+2   2.684863E+2   
4.254802E+3   7.003341E+1   7.003341E+1   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   -4.147209E-2   4.669164E-2   -5.604976E-5   1.483752E-7   -1.483752E-7   -5.604976E-5   5.604995E-5   1.798483E+2   2.698483E+2   
4.276565E+3   7.004241E+1   7.004241E+1   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   -4.336931E-2   4.758440E-2   -5.780416E-5   9.679515E-7   -9.679515E-7   -5.780416E-5   5.781226E-5   1.790407E+2   2.690407E+2   
4.298672E+3   7.003851E+1   7.003851E+1   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   -4.288306E-2   4.866712E-2   -5.820870E-5   -9.954528E-8   9.954528E-8   -5.820870E-5   5.820878E-5   -1.799020E+2   -8.990202E+1   
4.320491E+3   7.003619E+1   7.003619E+1   -1.499000E+3   -1.499000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   -4.449711E-2   5.098742E-2   -6.071776E-5   -4.226938E-7   4.226938E-7   -6.071776E-5   6.071923E-5   -1.796011E+2   -8.960114E+1   
4.342571E+3   7.005361E+1   7.005361E+1   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   -4.492202E-2   5.083096E-2   -6.087855E-5   -6.126212E-9   6.126212E-9   -6.087855E-5   6.087856E-5   -1.799942E+2   -8.999423E+1   
4.364647E+3   7.004760E+1   7.004760E+1   -1.399000E+3   -1.399000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   -4.603325E-2   5.417686E-2   -6.374472E-5   -1.371676E-6   1.371676E-6   -6.374472E-5   6.375948E-5   -1.787673E+2   -8.876728E+1   
4.386715E+3   7.001422E+1   7.001422E+1   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   -4.797774E-2   5.571143E-2   -6.594635E-5   -9.367274E-7   9.367274E-7   -6.594635E-5   6.595300E-5   -1.791862E+2   -8.918620E+1   
4.408819E+3   7.000369E+1   7.000369E+1   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   -4.879998E-2   5.628422E-2   -6.682775E-5   -7.030561E-7   7.030561E-7   -6.682775E-5   6.683144E-5   -1.793972E+2   -8.939725E+1   
4.430942E+3   7.002651E+1   7.002651E+1   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   -5.021586E-2   5.843146E-2   -6.910158E-5   -1.059625E-6   1.059625E-6   -6.910158E-5   6.910971E-5   -1.791215E+2   -8.912148E+1   
4.452957E+3   7.005010E+1   7.005010E+1   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   -4.934176E-2   5.916929E-2   -6.904171E-5   -2.188512E-6   2.188512E-6   -6.904171E-5   6.907639E-5   -1.781844E+2   -8.818442E+1   
4.475071E+3   7.002941E+1   7.002941E+1   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   -5.053245E-2   6.101249E-2   -7.097831E-5   -2.512873E-6   2.512873E-6   -7.097831E-5   7.102278E-5   -1.779724E+2   -8.797238E+1   
4.497114E+3   7.003170E+1   7.003170E+1   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   -5.176731E-2   6.324932E-2   -7.319858E-5   -3.061908E-6   3.061908E-6   -7.319858E-5   7.326259E-5   -1.776047E+2   -8.760471E+1   
4.519225E+3   7.003610E+1   7.003610E+1   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   -5.152555E-2   6.433139E-2   -7.375386E-5   -3.948148E-6   3.948148E-6   -7.375386E-5   7.385946E-5   -1.769358E+2   -8.693580E+1   
4.541292E+3   7.001260E+1   7.001260E+1   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   -5.469043E-2   6.602028E-2   -7.681049E-5   -2.711452E-6   2.711452E-6   -7.681049E-5   7.685833E-5   -1.779783E+2   -8.797827E+1   
4.563220E+3   7.003250E+1   7.003250E+1   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   -5.428515E-2   6.686886E-2   -7.711260E-5   -3.565985E-6   3.565985E-6   -7.711260E-5   7.719501E-5   -1.773523E+2   -8.735231E+1   
4.584897E+3   7.001019E+1   7.001019E+1   -9.000000E+2   -9.000000E+2   9.000000E+1   -8.990000E+2   -8.990000E+2   -5.521597E-2   6.803039E-2   -7.844457E-5   -3.636897E-6   3.636897E-6   -7.844457E-5   7.852883E-5   -1.773455E+2   -8.734552E+1   
4.606847E+3   7.003021E+1   7.003021E+1   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.490000E+2   -8.490000E+2   -5.682602E-2   6.982326E-2   -8.060765E-5   -3.618188E-6   3.618188E-6   -8.060765E-5   8.068882E-5   -1.774299E+2   -8.742992E+1   
4.628516E+3   7.000701E+1   7.000701E+1   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   -5.728682E-2   7.158917E-2   -8.204265E-5   -4.431866E-6   4.431866E-6   -8.204265E-5   8.216227E-5   -1.769079E+2   -8.690794E+1   
4.650238E+3   7.003439E+1   7.003439E+1   -7.500000E+2   -7.500000E+2   9.000000E+1   -7.490000E+2   -7.490000E+2   -5.795196E-2   7.365665E-2   -8.380041E-5   -5.291570E-6   5.291570E-6   -8.380041E-5   8.396731E-5   -1.763869E+2   -8.638686E+1   
4.672174E+3   7.002471E+1   7.002471E+1   -7.010000E+2   -7.010000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   -5.982061E-2   7.401559E-2   -8.518947E-5   -4.144116E-6   4.144116E-6   -8.518947E-5   8.529021E-5   -1.772150E+2   -8.721499E+1   
4.694142E+3   7.005609E+1   7.005609E+1   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.490000E+2   -6.490000E+2   -5.896098E-2   7.612785E-2   -8.603370E-5   -6.160861E-6   6.160861E-6   -8.603370E-5   8.625400E-5   -1.759040E+2   -8.590405E+1   
4.715755E+3   7.004830E+1   7.004830E+1   -6.000000E+2   -6.000000E+2   9.000000E+1   -6.000000E+2   -6.000000E+2   -6.011421E-2   7.705899E-2   -8.735312E-5   -5.916650E-6   5.916650E-6   -8.735312E-5   8.755327E-5   -1.761251E+2   -8.612513E+1   
4.737645E+3   7.003860E+1   7.003860E+1   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   -6.014459E-2   7.868927E-2   -8.843368E-5   -6.960014E-6   6.960014E-6   -8.843368E-5   8.870715E-5   -1.754999E+2   -8.549992E+1   
4.759257E+3   7.002111E+1   7.002111E+1   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   -6.272685E-2   8.007536E-2   -9.093290E-5   -5.956284E-6   5.956284E-6   -9.093290E-5   9.112777E-5   -1.762524E+2   -8.625237E+1   
4.780997E+3   7.003411E+1   7.003411E+1   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   -6.209212E-2   8.052543E-2   -9.083361E-5   -6.719992E-6   6.719992E-6   -9.083361E-5   9.108185E-5   -1.757689E+2   -8.576889E+1   
4.802627E+3   7.000201E+1   7.000201E+1   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   -6.260967E-2   8.236680E-2   -9.235285E-5   -7.541028E-6   7.541028E-6   -9.235285E-5   9.266022E-5   -1.753319E+2   -8.533190E+1   
4.824351E+3   6.999789E+1   6.999789E+1   -3.490000E+2   -3.490000E+2   9.000000E+1   -3.500000E+2   -3.500000E+2   -6.411940E-2   8.369121E-2   -9.414881E-5   -7.290249E-6   7.290249E-6   -9.414881E-5   9.443064E-5   -1.755722E+2   -8.557224E+1   
4.845934E+3   7.001000E+1   7.001000E+1   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   -6.535791E-2   8.590842E-2   -9.635856E-5   -7.823762E-6   7.823762E-6   -9.635856E-5   9.667566E-5   -1.753581E+2   -8.535809E+1   
4.867564E+3   7.002160E+1   7.002160E+1   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   -6.622399E-2   8.553075E-2   -9.664803E-5   -6.936268E-6   6.936268E-6   -9.664803E-5   9.689662E-5   -1.758950E+2   -8.589502E+1   
4.889167E+3   7.004641E+1   7.004641E+1   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   -6.757235E-2   8.766878E-2   -9.887414E-5   -7.336764E-6   7.336764E-6   -9.887414E-5   9.914597E-5   -1.757563E+2   -8.575625E+1   
4.910853E+3   7.002349E+1   7.002349E+1   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   -6.708548E-2   8.881036E-2   -9.931663E-5   -8.443197E-6   8.443197E-6   -9.931663E-5   9.967487E-5   -1.751408E+2   -8.514080E+1   
4.932475E+3   7.002871E+1   7.002871E+1   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   -6.998587E-2   9.010474E-2   -1.019528E-4   -7.144211E-6   7.144211E-6   -1.019528E-4   1.022028E-4   -1.759916E+2   -8.599162E+1   
4.954065E+3   7.001501E+1   7.001501E+1   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   -6.981867E-2   9.254040E-2   -1.034357E-4   -8.860246E-6   8.860246E-6   -1.034357E-4   1.038145E-4   -1.751040E+2   -8.510403E+1   
4.987154E+3   7.003661E+1   7.003661E+1   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   -7.031660E-2   9.180625E-2   -1.032654E-4   -8.011987E-6   8.011987E-6   -1.032654E-4   1.035758E-4   -1.755635E+2   -8.556352E+1   
5.009412E+3   7.000381E+1   7.000381E+1   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   -6.869766E-2   9.289049E-2   -1.029707E-4   -9.918254E-6   9.918254E-6   -1.029707E-4   1.034473E-4   -1.744982E+2   -8.449818E+1   
5.031619E+3   7.000359E+1   7.000359E+1   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   -6.936279E-2   9.238272E-2   -1.030512E-4   -9.094338E-6   9.094338E-6   -1.030512E-4   1.034517E-4   -1.749567E+2   -8.495668E+1   
5.053856E+3   7.001370E+1   7.001370E+1   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   -6.896427E-2   9.305832E-2   -1.032448E-4   -9.830785E-6   9.830785E-6   -1.032448E-4   1.037118E-4   -1.745608E+2   -8.456080E+1   
5.076079E+3   7.004110E+1   7.004110E+1   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   -6.900601E-2   9.230354E-2   -1.027791E-4   -9.306460E-6   9.306460E-6   -1.027791E-4   1.031995E-4   -1.748261E+2   -8.482608E+1   
5.098347E+3   7.004958E+1   7.004958E+1   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   -6.907993E-2   9.103277E-2   -1.019971E-4   -8.420994E-6   8.420994E-6   -1.019971E-4   1.023442E-4   -1.752803E+2   -8.528030E+1   
5.120614E+3   7.004989E+1   7.004989E+1   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   -6.915264E-2   9.204402E-2   -1.027007E-4   -9.028338E-6   9.028338E-6   -1.027007E-4   1.030968E-4   -1.749761E+2   -8.497609E+1   
5.142898E+3   7.000891E+1   7.000891E+1   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   -6.943334E-2   9.206519E-2   -1.028880E-4   -8.834562E-6   8.834562E-6   -1.028880E-4   1.032666E-4   -1.750923E+2   -8.509229E+1   
5.165174E+3   7.006921E+1   7.006921E+1   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   -7.014448E-2   9.349828E-2   -1.042610E-4   -9.245500E-6   9.245500E-6   -1.042610E-4   1.046702E-4   -1.749325E+2   -8.493247E+1   
5.187453E+3   7.000451E+1   7.000451E+1   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   -6.955055E-2   9.186086E-2   -1.028274E-4   -8.614289E-6   8.614289E-6   -1.028274E-4   1.031876E-4   -1.752113E+2   -8.521127E+1   
5.209674E+3   7.003021E+1   7.003021E+1   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   -7.064487E-2   9.271376E-2   -1.040595E-4   -8.362499E-6   8.362499E-6   -1.040595E-4   1.043949E-4   -1.754054E+2   -8.540543E+1   
5.231911E+3   7.001501E+1   7.001501E+1   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   -6.956435E-2   9.256593E-2   -1.032951E-4   -9.065037E-6   9.065037E-6   -1.032951E-4   1.036922E-4   -1.749847E+2   -8.498465E+1   
5.254163E+3   7.000259E+1   7.000259E+1   -2.300000E+1   -2.300000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   -7.029789E-2   9.214464E-2   -1.034743E-4   -8.247058E-6   8.247058E-6   -1.034743E-4   1.038024E-4   -1.754431E+2   -8.544307E+1   
5.275439E+3   7.001861E+1   7.001861E+1   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   -7.039484E-2   9.287269E-2   -1.040084E-4   -8.651328E-6   8.651328E-6   -1.040084E-4   1.043676E-4   -1.752451E+2   -8.524513E+1   
5.297723E+3   7.007849E+1   7.007849E+1   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   -6.989631E-2   9.303195E-2   -1.038039E-4   -9.124182E-6   9.124182E-6   -1.038039E-4   1.042041E-4   -1.749767E+2   -8.497671E+1   
5.319953E+3   6.997341E+1   6.997341E+1   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   -6.976714E-2   9.325961E-2   -1.038723E-4   -9.368553E-6   9.368553E-6   -1.038723E-4   1.042939E-4   -1.748463E+2   -8.484627E+1   
5.342136E+3   7.000640E+1   7.000640E+1   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   -7.058780E-2   9.279723E-2   -1.040785E-4   -8.459275E-6   8.459275E-6   -1.040785E-4   1.044217E-4   -1.753533E+2   -8.535334E+1   
5.364352E+3   7.001751E+1   7.001751E+1   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   -7.084920E-2   9.377225E-2   -1.048752E-4   -8.903382E-6   8.903382E-6   -1.048752E-4   1.052524E-4   -1.751475E+2   -8.514751E+1   
5.386624E+3   7.004440E+1   7.004440E+1   -1.100000E+1   -1.100000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   -7.011137E-2   9.278771E-2   -1.037778E-4   -8.805438E-6   8.805438E-6   -1.037778E-4   1.041507E-4   -1.751501E+2   -8.515013E+1   
5.407806E+3   7.003811E+1   7.003811E+1   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   -7.070255E-2   9.340840E-2   -1.045475E-4   -8.773970E-6   8.773970E-6   -1.045475E-4   1.049150E-4   -1.752028E+2   -8.520279E+1   
5.429898E+3   7.004958E+1   7.004958E+1   -7.000000E+0   -7.000000E+0   9.000000E+1   -6.000000E+0   -6.000000E+0   -6.931768E-2   9.352159E-2   -1.037651E-4   -9.872267E-6   9.872267E-6   -1.037651E-4   1.042336E-4   -1.745652E+2   -8.456521E+1   
5.450920E+3   6.999230E+1   6.999230E+1   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   -7.004142E-2   9.342711E-2   -1.041510E-4   -9.275200E-6   9.275200E-6   -1.041510E-4   1.045632E-4   -1.749109E+2   -8.491093E+1   
5.472942E+3   7.002670E+1   7.002670E+1   -3.000000E+0   -3.000000E+0   9.000000E+1   -2.000000E+0   -2.000000E+0   -7.030067E-2   9.348476E-2   -1.043488E-4   -9.121139E-6   9.121139E-6   -1.043488E-4   1.047467E-4   -1.750045E+2   -8.500447E+1   
5.493966E+3   7.004101E+1   7.004101E+1   -1.000000E+0   -1.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   -6.922442E-2   9.477003E-2   -1.045205E-4   -1.075744E-5   1.075744E-5   -1.045205E-4   1.050726E-4   -1.741237E+2   -8.412371E+1   
5.514929E+3   7.003079E+1   7.003079E+1   0.000000E+0   0.000000E+0   9.000000E+1   0.000000E+0   0.000000E+0   -7.048011E-2   9.378025E-2   -1.046522E-4   -9.181598E-6   9.181598E-6   -1.046522E-4   1.050542E-4   -1.749860E+2   -8.498603E+1   
5.536951E+3   7.002151E+1   7.002151E+1   1.000000E+0   1.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   -7.100875E-2   9.391402E-2   -1.050661E-4   -8.878056E-6   8.878056E-6   -1.050661E-4   1.054406E-4   -1.751700E+2   -8.517000E+1   
5.558667E+3   7.001980E+1   7.001980E+1   3.000000E+0   3.000000E+0   9.000000E+1   4.000000E+0   4.000000E+0   -7.003098E-2   9.409473E-2   -1.045793E-4   -9.719388E-6   9.719388E-6   -1.045793E-4   1.050300E-4   -1.746903E+2   -8.469030E+1   
5.580301E+3   7.003021E+1   7.003021E+1   5.000000E+0   5.000000E+0   9.000000E+1   6.000000E+0   6.000000E+0   -7.131002E-2   9.377530E-2   -1.051620E-4   -8.564542E-6   8.564542E-6   -1.051620E-4   1.055102E-4   -1.753440E+2   -8.534403E+1   
5.602031E+3   7.004260E+1   7.004260E+1   7.000000E+0   7.000000E+0   9.000000E+1   8.000000E+0   8.000000E+0   -7.113820E-2   9.381613E-2   -1.050824E-4   -8.718315E-6   8.718315E-6   -1.050824E-4   1.054435E-4   -1.752572E+2   -8.525723E+1   
5.623803E+3   7.005609E+1   7.005609E+1   9.000000E+0   9.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   -7.056479E-2   9.451970E-2   -1.051861E-4   -9.602396E-6   9.602396E-6   -1.051861E-4   1.056235E-4   -1.747840E+2   -8.478395E+1   
5.645804E+3   7.002120E+1   7.002120E+1   1.100000E+1   1.100000E+1   9.000000E+1   1.100000E+1   1.100000E+1   -7.050712E-2   9.348387E-2   -1.044759E-4   -8.967855E-6   8.967855E-6   -1.044759E-4   1.048600E-4   -1.750939E+2   -8.509395E+1   
5.667863E+3   7.006951E+1   7.006951E+1   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   -7.037183E-2   9.382412E-2   -1.046138E-4   -9.290367E-6   9.290367E-6   -1.046138E-4   1.050255E-4   -1.749251E+2   -8.492509E+1   
5.689772E+3   7.004641E+1   7.004641E+1   1.500000E+1   1.500000E+1   9.000000E+1   1.600000E+1   1.600000E+1   -7.029206E-2   9.467277E-2   -1.051172E-4   -9.904188E-6   9.904188E-6   -1.051172E-4   1.055828E-4   -1.746175E+2   -8.461746E+1   
5.711853E+3   7.002471E+1   7.002471E+1   1.700000E+1   1.700000E+1   9.000000E+1   1.800000E+1   1.800000E+1   -7.163794E-2   9.325868E-2   -1.050283E-4   -7.984244E-6   7.984244E-6   -1.050283E-4   1.053314E-4   -1.756527E+2   -8.565274E+1   
5.733997E+3   7.006710E+1   7.006710E+1   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   -7.042859E-2   9.449144E-2   -1.050835E-4   -9.684660E-6   9.684660E-6   -1.050835E-4   1.055289E-4   -1.747344E+2   -8.473441E+1   
5.755957E+3   7.000439E+1   7.000439E+1   2.100000E+1   2.100000E+1   9.000000E+1   2.100000E+1   2.100000E+1   -7.110477E-2   9.420550E-2   -1.053153E-4   -8.997600E-6   8.997600E-6   -1.053153E-4   1.056990E-4   -1.751168E+2   -8.511680E+1   
5.777991E+3   7.004421E+1   7.004421E+1   2.300000E+1   2.300000E+1   9.000000E+1   2.400000E+1   2.400000E+1   -7.020247E-2   9.320223E-2   -1.041041E-4   -9.009058E-6   9.009058E-6   -1.041041E-4   1.044932E-4   -1.750540E+2   -8.505401E+1   
5.800114E+3   7.002969E+1   7.002969E+1   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   -7.157322E-2   9.441380E-2   -1.057406E-4   -8.787303E-6   8.787303E-6   -1.057406E-4   1.061051E-4   -1.752495E+2   -8.524950E+1   
5.821957E+3   6.997921E+1   6.997921E+1   2.700000E+1   2.700000E+1   9.000000E+1   2.800000E+1   2.800000E+1   -7.121060E-2   9.369741E-2   -1.050499E-4   -8.587152E-6   8.587152E-6   -1.050499E-4   1.054002E-4   -1.753268E+2   -8.532683E+1   
5.844018E+3   7.002529E+1   7.002529E+1   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   -7.144192E-2   9.546155E-2   -1.063418E-4   -9.569403E-6   9.569403E-6   -1.063418E-4   1.067715E-4   -1.748580E+2   -8.485796E+1   
5.865983E+3   7.001190E+1   7.001190E+1   3.100000E+1   3.100000E+1   9.000000E+1   3.100000E+1   3.100000E+1   -7.036048E-2   9.442486E-2   -1.049981E-4   -9.691507E-6   9.691507E-6   -1.049981E-4   1.054444E-4   -1.747264E+2   -8.472644E+1   
5.888114E+3   7.001849E+1   7.001849E+1   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   -7.131277E-2   9.475866E-2   -1.058042E-4   -9.205398E-6   9.205398E-6   -1.058042E-4   1.062039E-4   -1.750276E+2   -8.502755E+1   
5.909964E+3   7.000491E+1   7.000491E+1   3.500000E+1   3.500000E+1   9.000000E+1   3.500000E+1   3.500000E+1   -7.125387E-2   9.604787E-2   -1.066074E-4   -1.009181E-5   1.009181E-5   -1.066074E-4   1.070840E-4   -1.745923E+2   -8.459231E+1   
5.932002E+3   7.003240E+1   7.003240E+1   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   -7.034422E-2   9.504093E-2   -1.053892E-4   -1.010630E-5   1.010630E-5   -1.053892E-4   1.058727E-4   -1.745224E+2   -8.452237E+1   
5.953977E+3   7.001891E+1   7.001891E+1   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   -7.158765E-2   9.371122E-2   -1.052920E-4   -8.317296E-6   8.317296E-6   -1.052920E-4   1.056199E-4   -1.754834E+2   -8.548343E+1   
5.975819E+3   7.003188E+1   7.003188E+1   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   -7.084489E-2   9.518391E-2   -1.057919E-4   -9.829473E-6   9.829473E-6   -1.057919E-4   1.062476E-4   -1.746917E+2   -8.469170E+1   
5.997695E+3   7.001321E+1   7.001321E+1   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   -7.204844E-2   9.572360E-2   -1.068875E-4   -9.292122E-6   9.292122E-6   -1.068875E-4   1.072906E-4   -1.750316E+2   -8.503156E+1   
6.019560E+3   6.999899E+1   6.999899E+1   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   -7.166743E-2   9.493725E-2   -1.061398E-4   -9.059834E-6   9.059834E-6   -1.061398E-4   1.065257E-4   -1.751212E+2   -8.512120E+1   
6.041435E+3   7.005120E+1   7.005120E+1   4.700000E+1   4.700000E+1   9.000000E+1   4.800000E+1   4.800000E+1   -7.153916E-2   9.558551E-2   -1.064827E-4   -9.578521E-6   9.578521E-6   -1.064827E-4   1.069126E-4   -1.748599E+2   -8.485986E+1   
6.063580E+3   7.002010E+1   7.002010E+1   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   -7.071727E-2   9.492587E-2   -1.055449E-4   -9.755164E-6   9.755164E-6   -1.055449E-4   1.059948E-4   -1.747193E+2   -8.471935E+1   
6.097089E+3   7.001989E+1   7.001989E+1   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   -7.199293E-2   9.718000E-2   -1.078017E-4   -1.028534E-5   1.028534E-5   -1.078017E-4   1.082913E-4   -1.745499E+2   -8.454992E+1   
6.119657E+3   7.001241E+1   7.001241E+1   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   -7.253532E-2   9.708518E-2   -1.080753E-4   -9.822170E-6   9.822170E-6   -1.080753E-4   1.085207E-4   -1.748071E+2   -8.480707E+1   
6.141986E+3   7.003881E+1   7.003881E+1   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   -7.435922E-2   9.999516E-2   -1.110981E-4   -1.037562E-5   1.037562E-5   -1.110981E-4   1.115816E-4   -1.746645E+2   -8.466454E+1   
6.164363E+3   7.001739E+1   7.001739E+1   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   -7.615825E-2   9.991661E-2   -1.121592E-4   -8.993649E-6   8.993649E-6   -1.121592E-4   1.125192E-4   -1.754155E+2   -8.541546E+1   
6.187249E+3   6.999200E+1   6.999200E+1   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   -7.497771E-2   1.022921E-1   -1.129765E-4   -1.141984E-5   1.141984E-5   -1.129765E-4   1.135522E-4   -1.742281E+2   -8.422806E+1   
6.209552E+3   7.001019E+1   7.001019E+1   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   -7.678501E-2   1.033110E-1   -1.147574E-4   -1.074921E-5   1.074921E-5   -1.147574E-4   1.152598E-4   -1.746488E+2   -8.464878E+1   
6.231934E+3   7.002239E+1   7.002239E+1   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   -7.677979E-2   1.047741E-1   -1.157071E-4   -1.170961E-5   1.170961E-5   -1.157071E-4   1.162981E-4   -1.742213E+2   -8.422132E+1   
6.254611E+3   7.000741E+1   7.000741E+1   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   -7.945656E-2   1.049695E-1   -1.174893E-4   -9.857545E-6   9.857545E-6   -1.174893E-4   1.179021E-4   -1.752040E+2   -8.520402E+1   
6.276815E+3   7.000109E+1   7.000109E+1   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   -7.936453E-2   1.072566E-1   -1.189220E-4   -1.142088E-5   1.142088E-5   -1.189220E-4   1.194691E-4   -1.745143E+2   -8.451432E+1   
6.299444E+3   7.001721E+1   7.001721E+1   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   -7.969156E-2   1.078168E-1   -1.194890E-4   -1.154524E-5   1.154524E-5   -1.194890E-4   1.200455E-4   -1.744811E+2   -8.448111E+1   
6.322774E+3   7.002520E+1   7.002520E+1   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   -8.011892E-2   1.107117E-1   -1.216386E-4   -1.312176E-5   1.312176E-5   -1.216386E-4   1.223443E-4   -1.738430E+2   -8.384303E+1   
6.345398E+3   7.003570E+1   7.003570E+1   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   -8.128903E-2   1.104077E-1   -1.221640E-4   -1.205754E-5   1.205754E-5   -1.221640E-4   1.227576E-4   -1.743632E+2   -8.436319E+1   
6.368028E+3   7.000771E+1   7.000771E+1   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   -8.290982E-2   1.122472E-1   -1.243641E-4   -1.206138E-5   1.206138E-5   -1.243641E-4   1.249477E-4   -1.744605E+2   -8.446053E+1   
6.391362E+3   7.001760E+1   7.001760E+1   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   -8.381270E-2   1.134769E-1   -1.257232E-4   -1.219749E-5   1.219749E-5   -1.257232E-4   1.263135E-4   -1.744586E+2   -8.445859E+1   
6.413998E+3   7.000991E+1   7.000991E+1   7.980000E+2   7.980000E+2   9.000000E+1   7.980000E+2   7.980000E+2   -8.411981E-2   1.153501E-1   -1.271331E-4   -1.319503E-5   1.319503E-5   -1.271331E-4   1.278160E-4   -1.740745E+2   -8.407454E+1   
6.436549E+3   7.000961E+1   7.000961E+1   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   -8.396919E-2   1.160582E-1   -1.275011E-4   -1.376935E-5   1.376935E-5   -1.275011E-4   1.282425E-4   -1.738363E+2   -8.383629E+1   
6.459893E+3   7.000689E+1   7.000689E+1   8.980000E+2   8.980000E+2   9.000000E+1   8.980000E+2   8.980000E+2   -8.525371E-2   1.175351E-1   -1.292572E-4   -1.378484E-5   1.378484E-5   -1.292572E-4   1.299902E-4   -1.739126E+2   -8.391261E+1   
6.482527E+3   7.001721E+1   7.001721E+1   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   -8.498191E-2   1.176928E-1   -1.291919E-4   -1.408896E-5   1.408896E-5   -1.291919E-4   1.299578E-4   -1.737762E+2   -8.377623E+1   
6.505071E+3   7.001580E+1   7.001580E+1   9.980000E+2   9.980000E+2   9.000000E+1   9.980000E+2   9.980000E+2   -8.837872E-2   1.206383E-1   -1.332103E-4   -1.350227E-5   1.350227E-5   -1.332103E-4   1.338929E-4   -1.742122E+2   -8.421224E+1   
6.528498E+3   6.997201E+1   6.997201E+1   1.048000E+3   1.048000E+3   9.000000E+1   1.048000E+3   1.048000E+3   -8.775837E-2   1.210190E-1   -1.330747E-4   -1.421001E-5   1.421001E-5   -1.330747E-4   1.338313E-4   -1.739049E+2   -8.390493E+1   
6.551288E+3   7.003381E+1   7.003381E+1   1.098000E+3   1.098000E+3   9.000000E+1   1.098000E+3   1.098000E+3   -8.863307E-2   1.233237E-1   -1.351165E-4   -1.506975E-5   1.506975E-5   -1.351165E-4   1.359543E-4   -1.736360E+2   -8.363601E+1   
6.574174E+3   7.002700E+1   7.002700E+1   1.148000E+3   1.148000E+3   9.000000E+1   1.149000E+3   1.149000E+3   -8.941078E-2   1.237968E-1   -1.359054E-4   -1.480383E-5   1.480383E-5   -1.359054E-4   1.367093E-4   -1.737834E+2   -8.378343E+1   
6.597448E+3   7.000689E+1   7.000689E+1   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   -8.937179E-2   1.250810E-1   -1.367177E-4   -1.567224E-5   1.567224E-5   -1.367177E-4   1.376131E-4   -1.734606E+2   -8.346061E+1   
6.620008E+3   7.001431E+1   7.001431E+1   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   -9.275154E-2   1.276412E-1   -1.404747E-4   -1.484626E-5   1.484626E-5   -1.404747E-4   1.412570E-4   -1.739670E+2   -8.396701E+1   
6.642555E+3   7.002700E+1   7.002700E+1   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   -9.134850E-2   1.272491E-1   -1.393519E-4   -1.562767E-5   1.562767E-5   -1.393519E-4   1.402254E-4   -1.736013E+2   -8.360128E+1   
6.665612E+3   6.999859E+1   6.999859E+1   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   -9.348327E-2   1.299182E-1   -1.424101E-4   -1.579370E-5   1.579370E-5   -1.424101E-4   1.432832E-4   -1.736716E+2   -8.367159E+1   
6.688184E+3   6.997299E+1   6.997299E+1   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   -9.328902E-2   1.310880E-1   -1.430518E-4   -1.670215E-5   1.670215E-5   -1.430518E-4   1.440236E-4   -1.733405E+2   -8.334053E+1   
6.710679E+3   6.999700E+1   6.999700E+1   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   -9.473292E-2   1.328170E-1   -1.450707E-4   -1.676462E-5   1.676462E-5   -1.450707E-4   1.460361E-4   -1.734080E+2   -8.340804E+1   
6.733468E+3   7.001199E+1   7.001199E+1   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   -9.455558E-2   1.338874E-1   -1.456582E-4   -1.759558E-5   1.759558E-5   -1.456582E-4   1.467171E-4   -1.731120E+2   -8.311201E+1   
6.756015E+3   6.998510E+1   6.998510E+1   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   -9.755029E-2   1.371582E-1   -1.496398E-4   -1.751890E-5   1.751890E-5   -1.496398E-4   1.506618E-4   -1.733226E+2   -8.332256E+1   
6.778586E+3   7.000771E+1   7.000771E+1   1.599000E+3   1.599000E+3   9.000000E+1   1.599000E+3   1.599000E+3   -9.609142E-2   1.367691E-1   -1.484845E-4   -1.834361E-5   1.834361E-5   -1.484845E-4   1.496133E-4   -1.729574E+2   -8.295743E+1   
6.801465E+3   7.000329E+1   7.000329E+1   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   -9.755118E-2   1.384580E-1   -1.504870E-4   -1.836808E-5   1.836808E-5   -1.504870E-4   1.516038E-4   -1.730410E+2   -8.304104E+1   
6.823965E+3   7.003240E+1   7.003240E+1   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   -9.940336E-2   1.388728E-1   -1.519022E-4   -1.726933E-5   1.726933E-5   -1.519022E-4   1.528807E-4   -1.735141E+2   -8.351405E+1   
6.846496E+3   7.000179E+1   7.000179E+1   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   -9.728884E-2   1.398536E-1   -1.512337E-4   -1.947451E-5   1.947451E-5   -1.512337E-4   1.524824E-4   -1.726623E+2   -8.266235E+1   
6.869287E+3   7.000030E+1   7.000030E+1   1.799000E+3   1.799000E+3   9.000000E+1   1.799000E+3   1.799000E+3   -1.015408E-1   1.426102E-1   -1.556578E-4   -1.813180E-5   1.813180E-5   -1.556578E-4   1.567102E-4   -1.733558E+2   -8.335584E+1   
6.891863E+3   7.002700E+1   7.002700E+1   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   -1.002768E-1   1.425378E-1   -1.548291E-4   -1.901935E-5   1.901935E-5   -1.548291E-4   1.559929E-4   -1.729968E+2   -8.299682E+1   
6.913906E+3   6.999639E+1   6.999639E+1   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   -1.023519E-1   1.454133E-1   -1.579849E-4   -1.936447E-5   1.936447E-5   -1.579849E-4   1.591673E-4   -1.730120E+2   -8.301202E+1   
6.936659E+3   7.001940E+1   7.001940E+1   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   -1.035441E-1   1.485887E-1   -1.607900E-4   -2.055861E-5   2.055861E-5   -1.607900E-4   1.620990E-4   -1.727137E+2   -8.271370E+1   
6.959238E+3   7.000530E+1   7.000530E+1   1.999000E+3   1.999000E+3   9.000000E+1   2.000000E+3   2.000000E+3   -1.027817E-1   1.465976E-1   -1.590219E-4   -1.982078E-5   1.982078E-5   -1.590219E-4   1.602524E-4   -1.728952E+2   -8.289519E+1   
6.997190E+3   7.003951E+1   7.003951E+1   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   -1.115591E-1   1.613411E-1   -1.740508E-4   -2.296769E-5   2.296769E-5   -1.740508E-4   1.755596E-4   -1.724827E+2   -8.248270E+1   
7.024099E+3   7.003460E+1   7.003460E+1   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   -1.202738E-1   1.746019E-1   -1.880753E-4   -2.519152E-5   2.519152E-5   -1.880753E-4   1.897549E-4   -1.723710E+2   -8.237099E+1   
7.050456E+3   7.000549E+1   7.000549E+1   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -1.312959E-1   1.923355E-1   -2.064393E-4   -2.863294E-5   2.863294E-5   -2.064393E-4   2.084156E-4   -1.721035E+2   -8.210351E+1   
7.076323E+3   7.003909E+1   7.003909E+1   3.998000E+3   3.998000E+3   9.000000E+1   4.000000E+3   4.000000E+3   -1.385970E-1   2.068465E-1   -2.204041E-4   -3.271975E-5   3.271975E-5   -2.204041E-4   2.228195E-4   -1.715559E+2   -8.155592E+1   
7.102936E+3   7.003811E+1   7.003811E+1   4.498000E+3   4.498000E+3   9.000000E+1   4.499000E+3   4.499000E+3   -1.468632E-1   2.194661E-1   -2.337337E-4   -3.485613E-5   3.485613E-5   -2.337337E-4   2.363184E-4   -1.715181E+2   -8.151813E+1   
7.128843E+3   7.000170E+1   7.000170E+1   4.998000E+3   4.998000E+3   9.000000E+1   4.999000E+3   4.999000E+3   -1.482493E-1   2.244052E-1   -2.378074E-4   -3.705996E-5   3.705996E-5   -2.378074E-4   2.406778E-4   -1.711423E+2   -8.114226E+1   
7.154514E+3   7.001669E+1   7.001669E+1   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -1.415876E-1   2.210338E-1   -2.314931E-4   -3.978305E-5   3.978305E-5   -2.314931E-4   2.348866E-4   -1.702487E+2   -8.024873E+1   
7.180913E+3   6.999569E+1   6.999569E+1   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -1.252724E-1   2.072144E-1   -2.124058E-4   -4.281553E-5   4.281553E-5   -2.124058E-4   2.166781E-4   -1.686034E+2   -7.860337E+1   
7.206591E+3   7.002331E+1   7.002331E+1   6.498000E+3   6.498000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -1.089023E-1   1.898064E-1   -1.909474E-4   -4.354257E-5   4.354257E-5   -1.909474E-4   1.958491E-4   -1.671542E+2   -7.715424E+1   
7.232768E+3   7.001669E+1   7.001669E+1   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -8.960903E-2   1.705832E-1   -1.664995E-4   -4.524486E-5   4.524486E-5   -1.664995E-4   1.725375E-4   -1.647975E+2   -7.479745E+1   
7.258461E+3   7.001281E+1   7.001281E+1   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -7.511791E-2   1.563928E-1   -1.482984E-4   -4.668566E-5   4.668566E-5   -1.482984E-4   1.554734E-4   -1.625255E+2   -7.252553E+1   
7.283837E+3   7.005209E+1   7.005209E+1   7.999000E+3   7.999000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -7.015707E-2   1.532939E-1   -1.432131E-4   -4.832889E-5   4.832889E-5   -1.432131E-4   1.511478E-4   -1.613524E+2   -7.135245E+1   
7.310275E+3   6.997070E+1   6.997070E+1   8.498000E+3   8.498000E+3   9.000000E+1   8.499000E+3   8.499000E+3   -7.158826E-2   1.587689E-1   -1.476637E-4   -5.084975E-5   5.084975E-5   -1.476637E-4   1.561739E-4   -1.609982E+2   -7.099825E+1   
7.336681E+3   7.005529E+1   7.005529E+1   8.998000E+3   8.998000E+3   9.000000E+1   8.999000E+3   8.999000E+3   -7.384167E-2   1.661090E-1   -1.538374E-4   -5.398176E-5   5.398176E-5   -1.538374E-4   1.630336E-4   -1.606640E+2   -7.066395E+1   
7.363108E+3   6.998681E+1   6.998681E+1   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -8.083346E-2   1.798790E-1   -1.671283E-4   -5.781291E-5   5.781291E-5   -1.671283E-4   1.768452E-4   -1.609185E+2   -7.091851E+1   
7.388558E+3   6.997909E+1   6.997909E+1   9.999000E+3   9.999000E+3   9.000000E+1   1.000000E+4   1.000000E+4   -8.800111E-2   1.921694E-1   -1.795643E-4   -6.054656E-5   6.054656E-5   -1.795643E-4   1.894973E-4   -1.613666E+2   -7.136661E+1   
@@END Data.
@Time at end of measurement: 17:29:14
@NO Instrument  Changes.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -9499.000      -9998.000      249.500        Coercive Field: Field at which M//H changes sign
Ms  emu                                 2.822E-4       -2.400E-4      2.611E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -1.047E-4      1.387E-4       1.217E-4       Remanent Magnetization: M at H=0        
S                                       0.371          0.578          0.474          Squareness: Mr/Ms                       
S*                                      1.393          1.411          1.402          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
