@Filename: c:\vsm-lv\Will\data\AJA335e-FePtFeRh_1030nm_Tann_6\AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_80deg.VHD
@Measurement Controlfilename: C:\vsm-lv\Will\Recipes\10kOe OoP loop 80deg.VHC
@Signal Manipulation filename: c:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA335e-FePtFeRh_1030nm_Tann_6
@Date: 07 November 2019    (2019-07-11)
@Time: 10:49:22
@Test ID: AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_80deg
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 90.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Sample Temperature to 80.1216 [degC] and wait 60.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Applied Field to 9999.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 3:      Set Auto Range Signal to 13.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 5
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 5.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 10000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To: 50.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: 50.0000 [Oe] To: -50.0000 [Oe] Min Stepsize/Sweeprate =  2.0000 [Oe] Max Stepsize/Sweeprate =  2.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -50.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -10000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 4 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 50 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.706
@Y Coils Correction Factor: 0.964
@Sample Shape Correction Factor: 0.919
@Coil Angle Alpha: 42.300
@Coil Angle Beta: -47.320
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
15000.000000   1.000000
15249.000000   1.000524
15499.000000   1.000702
15750.000000   1.001233
16000.000000   1.001406
16250.000000   1.001585
16499.000000   1.001758
16749.000000   1.001937
16999.000000   1.002110
17249.000000   1.001937
17499.000000   1.002289
17749.000000   1.002289
17999.000000   1.002289
18249.000000   1.002462
18499.000000   1.002462
18748.000000   1.002462
18999.000000   1.002462
19249.000000   1.002462
19499.000000   1.002642
19749.000000   1.002642
19999.000000   1.002462
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = No
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 25 October 2019  12:02:56
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 5
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 10:49:22
@@Data
New Section: Section 0: 
2.967700E+1   8.007339E+1   8.007339E+1   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -2.763100E-1   3.491270E-1   -3.982105E-4   -2.388194E-5   2.388194E-5   -3.982105E-4   3.989260E-4   -1.765679E+2   -8.656790E+1   
5.464700E+1   8.001620E+1   8.001620E+1   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -2.535703E-1   3.199743E-1   -3.651649E-4   -2.164169E-5   2.164169E-5   -3.651649E-4   3.658057E-4   -1.766083E+2   -8.660830E+1   
7.976300E+1   8.007150E+1   8.007150E+1   8.998000E+3   8.998000E+3   9.000000E+1   8.998000E+3   8.998000E+3   -2.358206E-1   2.960987E-1   -3.386413E-4   -1.916075E-5   1.916075E-5   -3.386413E-4   3.391829E-4   -1.767616E+2   -8.676159E+1   
1.048620E+2   8.000411E+1   8.000411E+1   8.497000E+3   8.497000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -2.149814E-1   2.718049E-1   -3.099352E-4   -1.869141E-5   1.869141E-5   -3.099352E-4   3.104983E-4   -1.765488E+2   -8.654882E+1   
1.306170E+2   8.005001E+1   8.005001E+1   7.998000E+3   7.998000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -1.959614E-1   2.499527E-1   -2.839440E-4   -1.847285E-5   1.847285E-5   -2.839440E-4   2.845443E-4   -1.762777E+2   -8.627769E+1   
1.564640E+2   8.004070E+1   8.004070E+1   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -1.757192E-1   2.252154E-1   -2.553182E-4   -1.727208E-5   1.727208E-5   -2.553182E-4   2.559018E-4   -1.761299E+2   -8.612988E+1   
1.813650E+2   8.005490E+1   8.005490E+1   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -1.544020E-1   1.980084E-1   -2.244194E-4   -1.525176E-5   1.525176E-5   -2.244194E-4   2.249370E-4   -1.761121E+2   -8.611210E+1   
2.066860E+2   8.004110E+1   8.004110E+1   6.498000E+3   6.498000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -1.353245E-1   1.749431E-1   -1.976025E-4   -1.428264E-5   1.428264E-5   -1.976025E-4   1.981180E-4   -1.758659E+2   -8.586587E+1   
2.320120E+2   8.004720E+1   8.004720E+1   5.998000E+3   5.998000E+3   9.000000E+1   5.998000E+3   5.998000E+3   -1.164230E-1   1.511488E-1   -1.704198E-4   -1.270678E-5   1.270678E-5   -1.704198E-4   1.708928E-4   -1.757358E+2   -8.573582E+1   
2.574660E+2   8.002670E+1   8.002670E+1   5.498000E+3   5.498000E+3   9.000000E+1   5.498000E+3   5.498000E+3   -9.232049E-2   1.212322E-1   -1.360341E-4   -1.097512E-5   1.097512E-5   -1.360341E-4   1.364761E-4   -1.753874E+2   -8.538742E+1   
2.829830E+2   8.003579E+1   8.003579E+1   4.998000E+3   4.998000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -7.845705E-2   1.020436E-1   -1.149657E-4   -8.683959E-6   8.683959E-6   -1.149657E-4   1.152932E-4   -1.756804E+2   -8.568035E+1   
3.085620E+2   8.002081E+1   8.002081E+1   4.498000E+3   4.498000E+3   9.000000E+1   4.498000E+3   4.498000E+3   -5.999364E-2   7.962653E-2   -8.895079E-5   -7.684412E-6   7.684412E-6   -8.895079E-5   8.928210E-5   -1.750625E+2   -8.506251E+1   
3.348120E+2   7.998889E+1   7.998889E+1   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -4.112755E-2   5.612010E-2   -6.197740E-5   -6.270520E-6   6.270520E-6   -6.197740E-5   6.229380E-5   -1.742228E+2   -8.422280E+1   
3.606150E+2   8.006451E+1   8.006451E+1   3.498000E+3   3.498000E+3   9.000000E+1   3.498000E+3   3.498000E+3   -2.237634E-2   3.208025E-2   -3.472763E-5   -4.422925E-6   4.422925E-6   -3.472763E-5   3.500815E-5   -1.727419E+2   -8.274186E+1   
3.859780E+2   7.999520E+1   7.999520E+1   2.998000E+3   2.998000E+3   9.000000E+1   2.998000E+3   2.998000E+3   -5.514932E-3   1.100717E-2   -1.057844E-5   -3.117160E-6   3.117160E-6   -1.057844E-5   1.102815E-5   -1.635813E+2   -7.358128E+1   
4.118120E+2   8.003951E+1   8.003951E+1   2.498000E+3   2.498000E+3   9.000000E+1   2.498000E+3   2.498000E+3   1.020337E-2   -1.180115E-2   1.399416E-5   1.685325E-7   -1.685325E-7   1.399416E-5   1.399518E-5   6.899830E-1   9.068998E+1   
4.376680E+2   8.004571E+1   8.004571E+1   1.999000E+3   1.999000E+3   9.000000E+1   1.999000E+3   1.999000E+3   2.913565E-2   -3.552799E-2   4.115203E-5   1.677568E-6   -1.677568E-6   4.115203E-5   4.118621E-5   2.334377E+0   9.233438E+1   
4.715640E+2   8.002010E+1   8.002010E+1   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   3.085799E-2   -3.747120E-2   4.348245E-5   1.674085E-6   -1.674085E-6   4.348245E-5   4.351466E-5   2.204813E+0   9.220481E+1   
4.938430E+2   8.004131E+1   8.004131E+1   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   3.368845E-2   -4.004950E-2   4.691159E-5   1.266205E-6   -1.266205E-6   4.691159E-5   4.692868E-5   1.546112E+0   9.154611E+1   
5.161280E+2   8.000659E+1   8.000659E+1   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   3.439593E-2   -4.142761E-2   4.824654E-5   1.643899E-6   -1.643899E-6   4.824654E-5   4.827453E-5   1.951478E+0   9.195148E+1   
5.383590E+2   8.002010E+1   8.002010E+1   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   3.584399E-2   -4.443604E-2   5.110115E-5   2.539701E-6   -2.539701E-6   5.110115E-5   5.116422E-5   2.845230E+0   9.284523E+1   
5.606020E+2   8.003839E+1   8.003839E+1   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   3.977890E-2   -4.717760E-2   5.531944E-5   1.421670E-6   -1.421670E-6   5.531944E-5   5.533771E-5   1.472136E+0   9.147214E+1   
5.828770E+2   8.003149E+1   8.003149E+1   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   4.081220E-2   -4.936265E-2   5.738138E-5   2.085935E-6   -2.085935E-6   5.738138E-5   5.741929E-5   2.081907E+0   9.208191E+1   
6.051570E+2   8.003851E+1   8.003851E+1   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   4.355309E-2   -5.122120E-2   6.028638E-5   1.273753E-6   -1.273753E-6   6.028638E-5   6.029984E-5   1.210386E+0   9.121039E+1   
6.274230E+2   8.002319E+1   8.002319E+1   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   4.358623E-2   -5.184277E-2   6.071169E-5   1.655603E-6   -1.655603E-6   6.071169E-5   6.073426E-5   1.562065E+0   9.156206E+1   
6.494330E+2   8.004461E+1   8.004461E+1   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   4.660817E-2   -5.502422E-2   6.465204E-5   1.500427E-6   -1.500427E-6   6.465204E-5   6.466945E-5   1.329466E+0   9.132947E+1   
6.716610E+2   8.006631E+1   8.006631E+1   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   4.886009E-2   -5.803447E-2   6.800483E-5   1.802852E-6   -1.802852E-6   6.800483E-5   6.802872E-5   1.518593E+0   9.151859E+1   
6.939780E+2   8.005230E+1   8.005230E+1   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   5.031740E-2   -5.972795E-2   7.000875E-5   1.832136E-6   -1.832136E-6   7.000875E-5   7.003272E-5   1.499094E+0   9.149909E+1   
7.161800E+2   8.003939E+1   8.003939E+1   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   5.189065E-2   -6.188839E-2   7.238847E-5   2.080944E-6   -2.080944E-6   7.238847E-5   7.241838E-5   1.646623E+0   9.164662E+1   
7.384770E+2   8.002450E+1   8.002450E+1   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   5.339454E-2   -6.376166E-2   7.453830E-5   2.193310E-6   -2.193310E-6   7.453830E-5   7.457056E-5   1.685457E+0   9.168546E+1   
7.605020E+2   8.002068E+1   8.002068E+1   1.298000E+3   1.298000E+3   9.000000E+1   1.298000E+3   1.298000E+3   5.657843E-2   -6.632279E-2   7.817476E-5   1.512806E-6   -1.512806E-6   7.817476E-5   7.818940E-5   1.108626E+0   9.110863E+1   
7.827450E+2   8.005920E+1   8.005920E+1   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   5.766938E-2   -6.890902E-2   8.053363E-5   2.396706E-6   -2.396706E-6   8.053363E-5   8.056928E-5   1.704637E+0   9.170464E+1   
8.050360E+2   8.002529E+1   8.002529E+1   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   5.929170E-2   -7.103939E-2   8.292411E-5   2.589563E-6   -2.589563E-6   8.292411E-5   8.296453E-5   1.788657E+0   9.178866E+1   
8.272690E+2   8.003381E+1   8.003381E+1   1.148000E+3   1.148000E+3   9.000000E+1   1.149000E+3   1.149000E+3   6.026240E-2   -7.333052E-2   8.501642E-5   3.369482E-6   -3.369482E-6   8.501642E-5   8.508317E-5   2.269633E+0   9.226963E+1   
8.495560E+2   8.004571E+1   8.004571E+1   1.098000E+3   1.098000E+3   9.000000E+1   1.099000E+3   1.099000E+3   6.240810E-2   -7.494364E-2   8.739361E-5   2.837063E-6   -2.837063E-6   8.739361E-5   8.743965E-5   1.859343E+0   9.185934E+1   
8.718400E+2   8.002371E+1   8.002371E+1   1.048000E+3   1.048000E+3   9.000000E+1   1.048000E+3   1.048000E+3   6.448938E-2   -7.708323E-2   9.007385E-5   2.696487E-6   -2.696487E-6   9.007385E-5   9.011420E-5   1.714718E+0   9.171472E+1   
8.940270E+2   7.999560E+1   7.999560E+1   9.980000E+2   9.980000E+2   9.000000E+1   9.990000E+2   9.990000E+2   6.374879E-2   -7.946209E-2   9.116530E-5   4.799486E-6   -4.799486E-6   9.116530E-5   9.129155E-5   3.013610E+0   9.301361E+1   
9.158850E+2   8.002291E+1   8.002291E+1   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   6.891885E-2   -8.149612E-2   9.568642E-5   2.305337E-6   -2.305337E-6   9.568642E-5   9.571419E-5   1.380139E+0   9.138014E+1   
9.377300E+2   8.000491E+1   8.000491E+1   8.980000E+2   8.980000E+2   9.000000E+1   8.990000E+2   8.990000E+2   6.977296E-2   -8.285705E-2   9.710083E-5   2.563350E-6   -2.563350E-6   9.710083E-5   9.713466E-5   1.512192E+0   9.151219E+1   
9.595460E+2   8.006909E+1   8.006909E+1   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   6.963920E-2   -8.691039E-2   9.965803E-5   5.312239E-6   -5.312239E-6   9.965803E-5   9.979951E-5   3.051245E+0   9.305125E+1   
9.813980E+2   8.001141E+1   8.001141E+1   7.980000E+2   7.980000E+2   9.000000E+1   7.990000E+2   7.990000E+2   7.314400E-2   -8.831305E-2   1.027384E-4   3.637001E-6   -3.637001E-6   1.027384E-4   1.028028E-4   2.027458E+0   9.202746E+1   
1.003299E+3   7.999590E+1   7.999590E+1   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   7.447364E-2   -8.991820E-2   1.046059E-4   3.702958E-6   -3.702958E-6   1.046059E-4   1.046714E-4   2.027375E+0   9.202737E+1   
1.025187E+3   8.000079E+1   8.000079E+1   6.980000E+2   6.980000E+2   9.000000E+1   6.980000E+2   6.980000E+2   7.528236E-2   -9.135711E-2   1.060430E-4   4.045521E-6   -4.045521E-6   1.060430E-4   1.061201E-4   2.184764E+0   9.218476E+1   
1.047009E+3   8.005319E+1   8.005319E+1   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   7.658253E-2   -9.373177E-2   1.083934E-4   4.636367E-6   -4.636367E-6   1.083934E-4   1.084925E-4   2.449249E+0   9.244925E+1   
1.068875E+3   7.999459E+1   7.999459E+1   5.980000E+2   5.980000E+2   9.000000E+1   5.990000E+2   5.990000E+2   7.841714E-2   -9.528357E-2   1.105383E-4   4.293953E-6   -4.293953E-6   1.105383E-4   1.106217E-4   2.224583E+0   9.222458E+1   
1.090743E+3   8.004391E+1   8.004391E+1   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   7.985233E-2   -9.774784E-2   1.130306E-4   4.843514E-6   -4.843514E-6   1.130306E-4   1.131343E-4   2.453701E+0   9.245370E+1   
1.112563E+3   8.005981E+1   8.005981E+1   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   8.124946E-2   -9.979665E-2   1.152287E-4   5.149607E-6   -5.149607E-6   1.152287E-4   1.153437E-4   2.558863E+0   9.255886E+1   
1.134424E+3   8.007009E+1   8.007009E+1   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   8.355285E-2   -1.011827E-1   1.175555E-4   4.352132E-6   -4.352132E-6   1.175555E-4   1.176361E-4   2.120232E+0   9.212023E+1   
1.156305E+3   8.001959E+1   8.001959E+1   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   8.542798E-2   -1.035475E-1   1.202550E-4   4.511238E-6   -4.511238E-6   1.202550E-4   1.203396E-4   2.148383E+0   9.214838E+1   
1.178142E+3   8.003149E+1   8.003149E+1   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   8.664288E-2   -1.056558E-1   1.223792E-4   4.990999E-6   -4.990999E-6   1.223792E-4   1.224809E-4   2.335404E+0   9.233540E+1   
1.200030E+3   8.005279E+1   8.005279E+1   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   8.678767E-2   -1.072542E-1   1.235097E-4   5.928893E-6   -5.928893E-6   1.235097E-4   1.236519E-4   2.748286E+0   9.274829E+1   
1.221940E+3   8.006460E+1   8.006460E+1   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   8.895920E-2   -1.087329E-1   1.258153E-4   5.289517E-6   -5.289517E-6   1.258153E-4   1.259265E-4   2.407407E+0   9.240741E+1   
1.243770E+3   8.004199E+1   8.004199E+1   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   8.967400E-2   -1.115763E-1   1.281091E-4   6.619734E-6   -6.619734E-6   1.281091E-4   1.282800E-4   2.957993E+0   9.295799E+1   
1.265605E+3   8.002151E+1   8.002151E+1   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   9.324951E-2   -1.129912E-1   1.312412E-4   4.900214E-6   -4.900214E-6   1.312412E-4   1.313326E-4   2.138287E+0   9.213829E+1   
1.287376E+3   8.002401E+1   8.002401E+1   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   9.352742E-2   -1.159155E-1   1.333176E-4   6.606521E-6   -6.606521E-6   1.333176E-4   1.334812E-4   2.836958E+0   9.283696E+1   
1.309151E+3   7.997119E+1   7.997119E+1   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   9.463259E-2   -1.176317E-1   1.351186E-4   6.911101E-6   -6.911101E-6   1.351186E-4   1.352952E-4   2.928036E+0   9.292804E+1   
1.342346E+3   8.000839E+1   8.000839E+1   4.600000E+1   4.600000E+1   9.000000E+1   4.700000E+1   4.700000E+1   9.603406E-2   -1.180944E-1   1.362864E-4   6.176992E-6   -6.176992E-6   1.362864E-4   1.364263E-4   2.595076E+0   9.259508E+1   
1.361321E+3   8.001040E+1   8.001040E+1   4.700000E+1   4.700000E+1   9.000000E+1   4.700000E+1   4.700000E+1   9.507805E-2   -1.172581E-1   1.351506E-4   6.337333E-6   -6.337333E-6   1.351506E-4   1.352991E-4   2.684683E+0   9.268468E+1   
1.383439E+3   8.002041E+1   8.002041E+1   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   9.458839E-2   -1.175532E-1   1.350401E-4   6.892440E-6   -6.892440E-6   1.350401E-4   1.352159E-4   2.921838E+0   9.292184E+1   
1.402532E+3   8.007641E+1   8.007641E+1   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   9.477247E-2   -1.180508E-1   1.354780E-4   7.081609E-6   -7.081609E-6   1.354780E-4   1.356630E-4   2.992201E+0   9.299220E+1   
1.424917E+3   8.000240E+1   8.000240E+1   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   9.501792E-2   -1.176017E-1   1.353372E-4   6.606451E-6   -6.606451E-6   1.353372E-4   1.354984E-4   2.794660E+0   9.279466E+1   
1.443931E+3   7.999511E+1   7.999511E+1   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   9.506333E-2   -1.182901E-1   1.358137E-4   7.022949E-6   -7.022949E-6   1.358137E-4   1.359952E-4   2.960138E+0   9.296014E+1   
1.466353E+3   8.008489E+1   8.008489E+1   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   9.602671E-2   -1.169175E-1   1.355153E-4   5.413038E-6   -5.413038E-6   1.355153E-4   1.356234E-4   2.287412E+0   9.228741E+1   
1.485386E+3   8.002029E+1   8.002029E+1   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   9.612611E-2   -1.171169E-1   1.357067E-4   5.469890E-6   -5.469890E-6   1.357067E-4   1.358169E-4   2.308155E+0   9.230816E+1   
1.507843E+3   8.001110E+1   8.001110E+1   3.000000E+1   3.000000E+1   9.000000E+1   3.100000E+1   3.100000E+1   9.625188E-2   -1.188988E-1   1.369449E-4   6.541787E-6   -6.541787E-6   1.369449E-4   1.371011E-4   2.734910E+0   9.273491E+1   
1.526901E+3   8.001061E+1   8.001061E+1   3.000000E+1   3.000000E+1   9.000000E+1   3.100000E+1   3.100000E+1   9.610588E-2   -1.172808E-1   1.358009E-4   5.591952E-6   -5.591952E-6   1.358009E-4   1.359160E-4   2.357970E+0   9.235797E+1   
1.549319E+3   8.004879E+1   8.004879E+1   2.600000E+1   2.600000E+1   9.000000E+1   2.700000E+1   2.700000E+1   9.433865E-2   -1.188270E-1   1.357153E-4   7.909927E-6   -7.909927E-6   1.357153E-4   1.359456E-4   3.335610E+0   9.333561E+1   
1.568319E+3   8.004901E+1   8.004901E+1   2.600000E+1   2.600000E+1   9.000000E+1   2.700000E+1   2.700000E+1   9.574628E-2   -1.191252E-1   1.367798E-4   7.063777E-6   -7.063777E-6   1.367798E-4   1.369621E-4   2.956324E+0   9.295632E+1   
1.590759E+3   7.998531E+1   7.998531E+1   2.300000E+1   2.300000E+1   9.000000E+1   2.300000E+1   2.300000E+1   9.626971E-2   -1.183281E-1   1.365843E-4   6.155527E-6   -6.155527E-6   1.365843E-4   1.367229E-4   2.580437E+0   9.258044E+1   
1.612189E+3   8.006109E+1   8.006109E+1   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   9.595308E-2   -1.191528E-1   1.369256E-4   6.928857E-6   -6.928857E-6   1.369256E-4   1.371008E-4   2.896871E+0   9.289687E+1   
1.631273E+3   7.996261E+1   7.996261E+1   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   9.587456E-2   -1.185546E-1   1.364875E-4   6.595825E-6   -6.595825E-6   1.364875E-4   1.366467E-4   2.766695E+0   9.276669E+1   
1.653689E+3   8.002279E+1   8.002279E+1   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   9.618196E-2   -1.184607E-1   1.366164E-4   6.307081E-6   -6.307081E-6   1.366164E-4   1.367619E-4   2.643261E+0   9.264326E+1   
1.672715E+3   8.006851E+1   8.006851E+1   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   9.662866E-2   -1.193062E-1   1.374432E-4   6.529476E-6   -6.529476E-6   1.374432E-4   1.375982E-4   2.719889E+0   9.271989E+1   
1.695138E+3   8.003530E+1   8.003530E+1   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   9.566285E-2   -1.184429E-1   1.362839E-4   6.679414E-6   -6.679414E-6   1.362839E-4   1.364475E-4   2.805881E+0   9.280588E+1   
1.714236E+3   8.007021E+1   8.007021E+1   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   9.675322E-2   -1.196296E-1   1.377308E-4   6.648742E-6   -6.648742E-6   1.377308E-4   1.378912E-4   2.763719E+0   9.276372E+1   
1.736317E+3   8.003301E+1   8.003301E+1   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   9.650654E-2   -1.199904E-1   1.378133E-4   7.067070E-6   -7.067070E-6   1.378133E-4   1.379944E-4   2.935558E+0   9.293556E+1   
1.755044E+3   8.002700E+1   8.002700E+1   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   9.557387E-2   -1.178330E-1   1.358316E-4   6.346480E-6   -6.346480E-6   1.358316E-4   1.359798E-4   2.675093E+0   9.267509E+1   
1.777042E+3   7.997030E+1   7.997030E+1   5.000000E+0   5.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   9.603900E-2   -1.193191E-1   1.370871E-4   6.974026E-6   -6.974026E-6   1.370871E-4   1.372643E-4   2.912296E+0   9.291230E+1   
1.798069E+3   8.004180E+1   8.004180E+1   3.000000E+0   3.000000E+0   9.000000E+1   3.000000E+0   3.000000E+0   9.642679E-2   -1.190522E-1   1.371530E-4   6.512708E-6   -6.512708E-6   1.371530E-4   1.373075E-4   2.718647E+0   9.271865E+1   
1.819127E+3   8.005831E+1   8.005831E+1   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   9.532598E-2   -1.196351E-1   1.368520E-4   7.707990E-6   -7.707990E-6   1.368520E-4   1.370689E-4   3.223695E+0   9.322369E+1   
1.837840E+3   8.005389E+1   8.005389E+1   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   9.834367E-2   -1.185625E-1   1.380192E-4   4.774810E-6   -4.774810E-6   1.380192E-4   1.381018E-4   1.981372E+0   9.198137E+1   
1.859852E+3   7.999011E+1   7.999011E+1   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   9.827003E-2   -1.189086E-1   1.381990E-4   5.055520E-6   -5.055520E-6   1.381990E-4   1.382915E-4   2.095028E+0   9.209503E+1   
1.881888E+3   8.002810E+1   8.002810E+1   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   9.703484E-2   -1.187331E-1   1.373211E-4   5.854376E-6   -5.854376E-6   1.373211E-4   1.374458E-4   2.441198E+0   9.244120E+1   
1.903880E+3   8.006280E+1   8.006280E+1   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   9.711341E-2   -1.189841E-1   1.375331E-4   5.960333E-6   -5.960333E-6   1.375331E-4   1.376622E-4   2.481499E+0   9.248150E+1   
1.925907E+3   8.003420E+1   8.003420E+1   -8.000000E+0   -8.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   9.754231E-2   -1.198621E-1   1.383701E-4   6.217138E-6   -6.217138E-6   1.383701E-4   1.385097E-4   2.572639E+0   9.257264E+1   
1.948059E+3   8.005761E+1   8.005761E+1   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   9.578557E-2   -1.196277E-1   1.371314E-4   7.363249E-6   -7.363249E-6   1.371314E-4   1.373289E-4   3.073537E+0   9.307354E+1   
1.970305E+3   8.003640E+1   8.003640E+1   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   9.748155E-2   -1.197290E-1   1.382459E-4   6.175044E-6   -6.175044E-6   1.382459E-4   1.383837E-4   2.557537E+0   9.255754E+1   
1.992596E+3   8.001330E+1   8.001330E+1   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   9.582048E-2   -1.207267E-1   1.378687E-4   8.055875E-6   -8.055875E-6   1.378687E-4   1.381039E-4   3.344076E+0   9.334408E+1   
2.014832E+3   8.003420E+1   8.003420E+1   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   9.719133E-2   -1.196670E-1   1.380261E-4   6.349165E-6   -6.349165E-6   1.380261E-4   1.381720E-4   2.633735E+0   9.263374E+1   
2.037070E+3   8.004019E+1   8.004019E+1   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   9.688270E-2   -1.206101E-1   1.384495E-4   7.194020E-6   -7.194020E-6   1.384495E-4   1.386363E-4   2.974490E+0   9.297449E+1   
2.059343E+3   8.004531E+1   8.004531E+1   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   9.678758E-2   -1.201505E-1   1.380914E-4   6.963914E-6   -6.963914E-6   1.380914E-4   1.382668E-4   2.886967E+0   9.288697E+1   
2.081585E+3   8.002981E+1   8.002981E+1   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   9.693850E-2   -1.206622E-1   1.385179E-4   7.186832E-6   -7.186832E-6   1.385179E-4   1.387043E-4   2.970057E+0   9.297006E+1   
2.103859E+3   8.003311E+1   8.003311E+1   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   9.569044E-2   -1.208831E-1   1.378902E-4   8.254353E-6   -8.254353E-6   1.378902E-4   1.381370E-4   3.425739E+0   9.342574E+1   
2.126116E+3   8.002639E+1   8.002639E+1   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   9.746562E-2   -1.215513E-1   1.394229E-4   7.378223E-6   -7.378223E-6   1.394229E-4   1.396180E-4   3.029252E+0   9.302925E+1   
2.148383E+3   8.002349E+1   8.002349E+1   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   9.681089E-2   -1.206764E-1   1.384482E-4   7.290455E-6   -7.290455E-6   1.384482E-4   1.386401E-4   3.014317E+0   9.301432E+1   
2.170656E+3   8.001870E+1   8.001870E+1   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   9.794300E-2   -1.202530E-1   1.388724E-4   6.176313E-6   -6.176313E-6   1.388724E-4   1.390097E-4   2.546536E+0   9.254654E+1   
2.192937E+3   8.002181E+1   8.002181E+1   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   9.699805E-2   -1.203714E-1   1.383653E-4   6.952646E-6   -6.952646E-6   1.383653E-4   1.385399E-4   2.876605E+0   9.287661E+1   
2.215194E+3   8.000829E+1   8.000829E+1   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   9.782581E-2   -1.212543E-1   1.394522E-4   6.917657E-6   -6.917657E-6   1.394522E-4   1.396236E-4   2.839884E+0   9.283988E+1   
2.237433E+3   8.005020E+1   8.005020E+1   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   9.774844E-2   -1.200940E-1   1.386486E-4   6.216312E-6   -6.216312E-6   1.386486E-4   1.387879E-4   2.567137E+0   9.256714E+1   
2.259665E+3   7.999529E+1   7.999529E+1   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   9.710480E-2   -1.212464E-1   1.390012E-4   7.445720E-6   -7.445720E-6   1.390012E-4   1.392005E-4   3.066168E+0   9.306617E+1   
2.281890E+3   8.001669E+1   8.001669E+1   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   9.635316E-2   -1.206131E-1   1.381241E-4   7.587671E-6   -7.587671E-6   1.381241E-4   1.383323E-4   3.144310E+0   9.314431E+1   
2.304138E+3   8.000460E+1   8.000460E+1   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   9.797675E-2   -1.217569E-1   1.398728E-4   7.134549E-6   -7.134549E-6   1.398728E-4   1.400546E-4   2.919979E+0   9.291998E+1   
2.326393E+3   8.001110E+1   8.001110E+1   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   9.736807E-2   -1.210838E-1   1.390581E-4   7.144703E-6   -7.144703E-6   1.390581E-4   1.392415E-4   2.941229E+0   9.294123E+1   
2.348659E+3   8.002920E+1   8.002920E+1   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   9.682258E-2   -1.220839E-1   1.393722E-4   8.202023E-6   -8.202023E-6   1.393722E-4   1.396133E-4   3.367959E+0   9.336796E+1   
2.370893E+3   8.004360E+1   8.004360E+1   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   9.671089E-2   -1.208500E-1   1.384995E-4   7.477921E-6   -7.477921E-6   1.384995E-4   1.387012E-4   3.090536E+0   9.309054E+1   
2.393149E+3   7.998599E+1   7.998599E+1   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   9.839093E-2   -1.207843E-1   1.394954E-4   6.192408E-6   -6.192408E-6   1.394954E-4   1.396328E-4   2.541775E+0   9.254178E+1   
2.426481E+3   8.002361E+1   8.002361E+1   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   9.971812E-2   -1.226116E-1   1.415060E-4   6.405377E-6   -6.405377E-6   1.415060E-4   1.416509E-4   2.591767E+0   9.259177E+1   
2.448176E+3   8.001699E+1   8.001699E+1   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   9.983836E-2   -1.253157E-1   1.433415E-4   8.084291E-6   -8.084291E-6   1.433415E-4   1.435693E-4   3.227994E+0   9.322799E+1   
2.469808E+3   8.004141E+1   8.004141E+1   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   1.018068E-1   -1.270748E-1   1.457042E-4   7.778478E-6   -7.778478E-6   1.457042E-4   1.459117E-4   3.055858E+0   9.305586E+1   
2.491561E+3   8.004949E+1   8.004949E+1   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   1.020976E-1   -1.296322E-1   1.475496E-4   9.235321E-6   -9.235321E-6   1.475496E-4   1.478384E-4   3.581545E+0   9.358154E+1   
2.513739E+3   8.005651E+1   8.005651E+1   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   1.041488E-1   -1.298089E-1   1.489329E-4   7.833727E-6   -7.833727E-6   1.489329E-4   1.491387E-4   3.010929E+0   9.301093E+1   
2.535412E+3   7.999621E+1   7.999621E+1   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   1.060288E-1   -1.326603E-1   1.519522E-4   8.307317E-6   -8.307317E-6   1.519522E-4   1.521791E-4   3.129279E+0   9.312928E+1   
2.557142E+3   7.999029E+1   7.999029E+1   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   1.061853E-1   -1.334905E-1   1.525896E-4   8.734364E-6   -8.734364E-6   1.525896E-4   1.528394E-4   3.276086E+0   9.327609E+1   
2.578851E+3   8.001669E+1   8.001669E+1   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   1.081457E-1   -1.341182E-1   1.542105E-4   7.694728E-6   -7.694728E-6   1.542105E-4   1.544023E-4   2.856551E+0   9.285655E+1   
2.600584E+3   8.002950E+1   8.002950E+1   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   1.095023E-1   -1.367639E-1   1.567724E-4   8.421063E-6   -8.421063E-6   1.567724E-4   1.569984E-4   3.074700E+0   9.307470E+1   
2.622319E+3   8.001251E+1   8.001251E+1   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   1.106123E-1   -1.387047E-1   1.587226E-4   8.868901E-6   -8.868901E-6   1.587226E-4   1.589702E-4   3.198175E+0   9.319818E+1   
2.644048E+3   8.001461E+1   8.001461E+1   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   1.121309E-1   -1.406436E-1   1.609243E-4   9.013308E-6   -9.013308E-6   1.609243E-4   1.611765E-4   3.205765E+0   9.320576E+1   
2.665782E+3   8.004669E+1   8.004669E+1   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.490000E+2   -6.490000E+2   1.124414E-1   -1.413321E-1   1.615646E-4   9.233759E-6   -9.233759E-6   1.615646E-4   1.618283E-4   3.271016E+0   9.327102E+1   
2.687408E+3   8.002621E+1   8.002621E+1   -7.010000E+2   -7.010000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   1.145614E-1   -1.433072E-1   1.641617E-4   8.957061E-6   -8.957061E-6   1.641617E-4   1.644058E-4   3.123101E+0   9.312310E+1   
2.709137E+3   8.003188E+1   8.003188E+1   -7.510000E+2   -7.510000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   1.142306E-1   -1.442938E-1   1.645998E-4   9.846718E-6   -9.846718E-6   1.645998E-4   1.648940E-4   3.423479E+0   9.342348E+1   
2.730826E+3   8.003521E+1   8.003521E+1   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   1.163340E-1   -1.466445E-1   1.674311E-4   9.827805E-6   -9.827805E-6   1.674311E-4   1.677193E-4   3.359270E+0   9.335927E+1   
2.752528E+3   7.997961E+1   7.997961E+1   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   1.166647E-1   -1.482858E-1   1.687046E-4   1.065624E-5   -1.065624E-5   1.687046E-4   1.690408E-4   3.614293E+0   9.361429E+1   
2.774251E+3   8.002499E+1   8.002499E+1   -9.000000E+2   -9.000000E+2   9.000000E+1   -9.000000E+2   -9.000000E+2   1.177815E-1   -1.501493E-1   1.706086E-4   1.104855E-5   -1.104855E-5   1.706086E-4   1.709660E-4   3.705277E+0   9.370528E+1   
2.795882E+3   8.002090E+1   8.002090E+1   -9.510000E+2   -9.510000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   1.204733E-1   -1.511016E-1   1.728931E-4   9.680177E-6   -9.680177E-6   1.728931E-4   1.731638E-4   3.204610E+0   9.320461E+1   
2.817607E+3   8.003619E+1   8.003619E+1   -1.000000E+3   -1.000000E+3   9.000000E+1   -1.000000E+3   -1.000000E+3   1.203542E-1   -1.533203E-1   1.742645E-4   1.121877E-5   -1.121877E-5   1.742645E-4   1.746252E-4   3.683494E+0   9.368349E+1   
2.839732E+3   8.000570E+1   8.000570E+1   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   1.227355E-1   -1.541904E-1   1.763034E-4   1.002628E-5   -1.002628E-5   1.763034E-4   1.765883E-4   3.254875E+0   9.325487E+1   
2.861591E+3   7.999151E+1   7.999151E+1   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   1.238032E-1   -1.571669E-1   1.789020E-4   1.118258E-5   -1.118258E-5   1.789020E-4   1.792512E-4   3.576719E+0   9.357672E+1   
2.883432E+3   8.007079E+1   8.007079E+1   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   1.240161E-1   -1.590119E-1   1.802353E-4   1.223135E-5   -1.223135E-5   1.802353E-4   1.806499E-4   3.882324E+0   9.388232E+1   
2.906050E+3   7.999529E+1   7.999529E+1   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   1.254194E-1   -1.603538E-1   1.819769E-4   1.207075E-5   -1.207075E-5   1.819769E-4   1.823768E-4   3.794940E+0   9.379494E+1   
2.927834E+3   8.004431E+1   8.004431E+1   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   1.278676E-1   -1.614522E-1   1.842058E-4   1.097804E-5   -1.097804E-5   1.842058E-4   1.845326E-4   3.410600E+0   9.341060E+1   
2.949952E+3   8.004391E+1   8.004391E+1   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   1.288904E-1   -1.647631E-1   1.869945E-4   1.238609E-5   -1.238609E-5   1.869945E-4   1.874043E-4   3.789606E+0   9.378961E+1   
2.972501E+3   8.001861E+1   8.001861E+1   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   1.285045E-1   -1.647858E-1   1.867707E-4   1.268638E-5   -1.268638E-5   1.867707E-4   1.872011E-4   3.885841E+0   9.388584E+1   
2.994569E+3   8.003689E+1   8.003689E+1   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   1.307760E-1   -1.679782E-1   1.902543E-4   1.309347E-5   -1.309347E-5   1.902543E-4   1.907043E-4   3.936938E+0   9.393694E+1   
3.016452E+3   8.002459E+1   8.002459E+1   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   1.329922E-1   -1.698699E-1   1.928565E-4   1.269098E-5   -1.269098E-5   1.928565E-4   1.932736E-4   3.764937E+0   9.376494E+1   
3.038817E+3   8.003570E+1   8.003570E+1   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   1.344765E-1   -1.707952E-1   1.943768E-4   1.219809E-5   -1.219809E-5   1.943768E-4   1.947591E-4   3.590881E+0   9.359088E+1   
3.060928E+3   7.998370E+1   7.998370E+1   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   1.350183E-1   -1.733311E-1   1.963634E-4   1.345529E-5   -1.345529E-5   1.963634E-4   1.968238E-4   3.919917E+0   9.391992E+1   
3.083045E+3   8.001660E+1   8.001660E+1   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   1.352606E-1   -1.745976E-1   1.973380E-4   1.410400E-5   -1.410400E-5   1.973380E-4   1.978414E-4   4.088052E+0   9.408805E+1   
3.105375E+3   8.001141E+1   8.001141E+1   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   1.384261E-1   -1.755112E-1   1.998901E-4   1.236003E-5   -1.236003E-5   1.998901E-4   2.002719E-4   3.538329E+0   9.353833E+1   
3.127499E+3   8.000860E+1   8.000860E+1   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.698000E+3   -1.698000E+3   1.373339E-1   -1.783392E-1   2.010567E-4   1.501670E-5   -1.501670E-5   2.010567E-4   2.016167E-4   4.271426E+0   9.427143E+1   
3.149647E+3   8.002871E+1   8.002871E+1   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.748000E+3   -1.748000E+3   1.402227E-1   -1.783202E-1   2.028303E-4   1.286766E-5   -1.286766E-5   2.028303E-4   2.032380E-4   3.630009E+0   9.363001E+1   
3.172839E+3   8.002941E+1   8.002941E+1   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.798000E+3   -1.798000E+3   1.413996E-1   -1.816152E-1   2.057039E-4   1.415136E-5   -1.415136E-5   2.057039E-4   2.061901E-4   3.935451E+0   9.393545E+1   
3.194943E+3   8.002780E+1   8.002780E+1   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.848000E+3   -1.848000E+3   1.418015E-1   -1.833749E-1   2.070984E-4   1.500457E-5   -1.500457E-5   2.070984E-4   2.076413E-4   4.143918E+0   9.414392E+1   
3.217324E+3   8.003509E+1   8.003509E+1   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   1.430047E-1   -1.842002E-1   2.083799E-4   1.465419E-5   -1.465419E-5   2.083799E-4   2.088945E-4   4.022669E+0   9.402267E+1   
3.240109E+3   8.002291E+1   8.002291E+1   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   1.437570E-1   -1.865400E-1   2.103688E-4   1.562747E-5   -1.562747E-5   2.103688E-4   2.109485E-4   4.248474E+0   9.424847E+1   
3.262421E+3   7.999191E+1   7.999191E+1   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   1.443153E-1   -1.866467E-1   2.107835E-4   1.528427E-5   -1.528427E-5   2.107835E-4   2.113370E-4   4.147355E+0   9.414736E+1   
3.299962E+3   8.001330E+1   8.001330E+1   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.561219E-1   -2.063906E-1   2.309419E-4   1.945973E-5   -1.945973E-5   2.309419E-4   2.317603E-4   4.816504E+0   9.481650E+1   
3.326112E+3   8.002801E+1   8.002801E+1   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.685660E-1   -2.240551E-1   2.501401E-4   2.180421E-5   -2.180421E-5   2.501401E-4   2.510886E-4   4.981765E+0   9.498177E+1   
3.351332E+3   8.001660E+1   8.001660E+1   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.813937E-1   -2.424615E-1   2.700586E-4   2.435006E-5   -2.435006E-5   2.700586E-4   2.711542E-4   5.152190E+0   9.515219E+1   
3.376992E+3   8.004391E+1   8.004391E+1   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   1.938531E-1   -2.615397E-1   2.901871E-4   2.760748E-5   -2.760748E-5   2.901871E-4   2.914974E-4   5.434582E+0   9.543458E+1   
3.402672E+3   8.003869E+1   8.003869E+1   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   2.047591E-1   -2.770081E-1   3.070041E-4   2.965388E-5   -2.965388E-5   3.070041E-4   3.084329E-4   5.517150E+0   9.551715E+1   
3.427407E+3   8.004199E+1   8.004199E+1   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   2.095168E-1   -2.878245E-1   3.169901E-4   3.320638E-5   -3.320638E-5   3.169901E-4   3.187247E-4   5.980222E+0   9.598022E+1   
3.452660E+3   8.006640E+1   8.006640E+1   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   2.101231E-1   -2.907089E-1   3.192435E-4   3.464371E-5   -3.464371E-5   3.192435E-4   3.211177E-4   6.193395E+0   9.619340E+1   
3.478359E+3   8.001129E+1   8.001129E+1   -5.999000E+3   -5.999000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   2.001443E-1   -2.777162E-1   3.046122E-4   3.353005E-5   -3.353005E-5   3.046122E-4   3.064520E-4   6.281519E+0   9.628152E+1   
3.503118E+3   8.001000E+1   8.001000E+1   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.858448E-1   -2.617078E-1   2.853454E-4   3.364057E-5   -3.364057E-5   2.853454E-4   2.873216E-4   6.723802E+0   9.672380E+1   
3.527788E+3   7.999990E+1   7.999990E+1   -7.000000E+3   -7.000000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.745565E-1   -2.492582E-1   2.702582E-4   3.385057E-5   -3.385057E-5   2.702582E-4   2.723699E-4   7.139272E+0   9.713927E+1   
3.552952E+3   8.004809E+1   8.004809E+1   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.688655E-1   -2.425971E-1   2.624014E-4   3.370498E-5   -3.370498E-5   2.624014E-4   2.645573E-4   7.319459E+0   9.731946E+1   
3.578159E+3   7.999679E+1   7.999679E+1   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.710603E-1   -2.439801E-1   2.646591E-4   3.298579E-5   -3.298579E-5   2.646591E-4   2.667067E-4   7.104426E+0   9.710443E+1   
3.603359E+3   7.999771E+1   7.999771E+1   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.500000E+3   -8.500000E+3   1.759082E-1   -2.508816E-1   2.721512E-4   3.391213E-5   -3.391213E-5   2.721512E-4   2.742559E-4   7.102882E+0   9.710288E+1   
3.628503E+3   8.000039E+1   8.000039E+1   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.876311E-1   -2.671704E-1   2.900076E-4   3.589069E-5   -3.589069E-5   2.900076E-4   2.922200E-4   7.054925E+0   9.705493E+1   
3.653751E+3   8.001159E+1   8.001159E+1   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.975788E-1   -2.815836E-1   3.055449E-4   3.795599E-5   -3.795599E-5   3.055449E-4   3.078934E-4   7.081231E+0   9.708123E+1   
3.678903E+3   7.999630E+1   7.999630E+1   -9.999000E+3   -9.999000E+3   9.000000E+1   -9.999000E+3   -9.999000E+3   2.108735E-1   -3.003218E-1   3.259682E-4   4.037333E-5   -4.037333E-5   3.259682E-4   3.284590E-4   7.060506E+0   9.706051E+1   
3.715484E+3   8.002441E+1   8.002441E+1   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.908133E-1   -2.707144E-1   2.942831E-4   3.585404E-5   -3.585404E-5   2.942831E-4   2.964592E-4   6.946406E+0   9.694641E+1   
3.739674E+3   7.999841E+1   7.999841E+1   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.662412E-1   -2.441924E-1   2.618180E-4   3.668894E-5   -3.668894E-5   2.618180E-4   2.643761E-4   7.976998E+0   9.797700E+1   
3.764308E+3   8.010290E+1   8.010290E+1   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.502591E-1   -2.233476E-1   2.383612E-4   3.488207E-5   -3.488207E-5   2.383612E-4   2.409000E-4   8.325637E+0   9.832564E+1   
3.788955E+3   8.001861E+1   8.001861E+1   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.349336E-1   -2.030484E-1   2.156655E-4   3.294622E-5   -3.294622E-5   2.156655E-4   2.181675E-4   8.685658E+0   9.868566E+1   
3.813684E+3   8.004559E+1   8.004559E+1   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.262808E-1   -1.896173E-1   2.015685E-4   3.056521E-5   -3.056521E-5   2.015685E-4   2.038727E-4   8.622466E+0   9.862247E+1   
3.838870E+3   8.003930E+1   8.003930E+1   -7.000000E+3   -7.000000E+3   9.000000E+1   -6.999000E+3   -6.999000E+3   1.057908E-1   -1.637132E-1   1.720295E-4   2.878494E-5   -2.878494E-5   1.720295E-4   1.744211E-4   9.499053E+0   9.949905E+1   
3.863993E+3   8.010421E+1   8.010421E+1   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   9.483627E-2   -1.478220E-1   1.549071E-4   2.649797E-5   -2.649797E-5   1.549071E-4   1.571571E-4   9.706906E+0   9.970691E+1   
3.888224E+3   8.000881E+1   8.000881E+1   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   8.226801E-2   -1.304268E-1   1.358076E-4   2.442142E-5   -2.442142E-5   1.358076E-4   1.379859E-4   1.019419E+1   1.001942E+2   
3.912971E+3   8.001000E+1   8.001000E+1   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   7.008650E-2   -1.116714E-1   1.160611E-4   2.116943E-5   -2.116943E-5   1.160611E-4   1.179760E-4   1.033706E+1   1.003371E+2   
3.938168E+3   8.000930E+1   8.000930E+1   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   5.550344E-2   -9.182225E-2   9.411768E-5   1.897873E-5   -1.897873E-5   9.411768E-5   9.601213E-5   1.140075E+1   1.014007E+2   
3.962391E+3   8.002880E+1   8.002880E+1   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   4.205164E-2   -7.238745E-2   7.314346E-5   1.622217E-5   -1.622217E-5   7.314346E-5   7.492079E-5   1.250497E+1   1.025050E+2   
3.987106E+3   7.999310E+1   7.999310E+1   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   3.165136E-2   -5.696315E-2   5.666784E-5   1.383057E-5   -1.383057E-5   5.666784E-5   5.833120E-5   1.371569E+1   1.037157E+2   
4.011812E+3   8.003170E+1   8.003170E+1   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.861504E-2   -3.731044E-2   3.580859E-5   1.062425E-5   -1.062425E-5   3.580859E-5   3.735143E-5   1.652539E+1   1.065254E+2   
4.036042E+3   7.997689E+1   7.997689E+1   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   6.113183E-3   -1.847269E-2   1.581052E-5   7.555420E-6   -7.555420E-6   1.581052E-5   1.752304E-5   2.554187E+1   1.155419E+2   
4.060745E+3   8.003280E+1   8.003280E+1   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   -7.134193E-3   -2.840922E-4   -4.225666E-6   5.462402E-6   -5.462402E-6   -4.225666E-6   6.906091E-6   1.277252E+2   2.177252E+2   
4.085408E+3   8.002068E+1   8.002068E+1   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   -2.115715E-2   2.014961E-2   -2.620357E-5   2.475234E-6   -2.475234E-6   -2.620357E-5   2.632021E-5   1.746038E+2   2.646038E+2   
4.119151E+3   8.000439E+1   8.000439E+1   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   -2.054293E-2   2.280892E-2   -2.755581E-5   2.823568E-7   -2.823568E-7   -2.755581E-5   2.755726E-5   1.794129E+2   2.694129E+2   
4.141178E+3   8.002679E+1   8.002679E+1   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.899000E+3   -1.899000E+3   -2.319550E-2   2.523815E-2   -3.077789E-5   6.561244E-7   -6.561244E-7   -3.077789E-5   3.078488E-5   1.787788E+2   2.687788E+2   
4.163263E+3   8.003851E+1   8.003851E+1   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.849000E+3   -1.849000E+3   -2.369556E-2   2.619474E-2   -3.171006E-5   4.005932E-7   -4.005932E-7   -3.171006E-5   3.171259E-5   1.792762E+2   2.692762E+2   
4.185044E+3   8.001739E+1   8.001739E+1   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.799000E+3   -1.799000E+3   -2.548174E-2   2.915530E-2   -3.474254E-5   -2.138217E-7   2.138217E-7   -3.474254E-5   3.474320E-5   -1.796474E+2   -8.964738E+1   
4.207130E+3   8.009420E+1   8.009420E+1   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   -2.704638E-2   2.924057E-2   -3.576541E-5   8.876801E-7   -8.876801E-7   -3.576541E-5   3.577642E-5   1.785782E+2   2.685782E+2   
4.229163E+3   8.004470E+1   8.004470E+1   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   -2.728753E-2   3.112980E-2   -3.714493E-5   -1.690774E-7   1.690774E-7   -3.714493E-5   3.714532E-5   -1.797392E+2   -8.973920E+1   
4.251040E+3   8.008550E+1   8.008550E+1   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   -2.854415E-2   3.338105E-2   -3.938806E-5   -7.114507E-7   7.114507E-7   -3.938806E-5   3.939448E-5   -1.789652E+2   -8.896520E+1   
4.272874E+3   8.004040E+1   8.004040E+1   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.599000E+3   -1.599000E+3   -3.041375E-2   3.701594E-2   -4.291129E-5   -1.705017E-6   1.705017E-6   -4.291129E-5   4.294515E-5   -1.777246E+2   -8.772463E+1   
4.294742E+3   8.004171E+1   8.004171E+1   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   -3.114944E-2   3.676436E-2   -4.320228E-5   -9.964112E-7   9.964112E-7   -4.320228E-5   4.321377E-5   -1.786788E+2   -8.867877E+1   
4.316544E+3   8.008441E+1   8.008441E+1   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   -3.288711E-2   3.839465E-2   -4.533838E-5   -7.770065E-7   7.770065E-7   -4.533838E-5   4.534503E-5   -1.790182E+2   -8.901816E+1   
4.338597E+3   7.999429E+1   7.999429E+1   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   -3.385840E-2   4.001514E-2   -4.699429E-5   -1.118041E-6   1.118041E-6   -4.699429E-5   4.700758E-5   -1.786371E+2   -8.863713E+1   
4.360688E+3   8.000259E+1   8.000259E+1   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   -3.571205E-2   4.269651E-2   -4.988665E-5   -1.500028E-6   1.500028E-6   -4.988665E-5   4.990919E-5   -1.782777E+2   -8.827771E+1   
4.382473E+3   8.004269E+1   8.004269E+1   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   -3.565377E-2   4.439555E-2   -5.095718E-5   -2.653917E-6   2.653917E-6   -5.095718E-5   5.102624E-5   -1.770187E+2   -8.701865E+1   
4.404517E+3   7.999459E+1   7.999459E+1   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   -3.739634E-2   4.596882E-2   -5.305917E-5   -2.393620E-6   2.393620E-6   -5.305917E-5   5.311314E-5   -1.774170E+2   -8.741701E+1   
4.426595E+3   8.000659E+1   8.000659E+1   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.250000E+3   -1.250000E+3   -3.940827E-2   4.773474E-2   -5.545317E-5   -2.060040E-6   2.060040E-6   -5.545317E-5   5.549142E-5   -1.778725E+2   -8.787249E+1   
4.448612E+3   8.000710E+1   8.000710E+1   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.200000E+3   -1.200000E+3   -3.944695E-2   4.960746E-2   -5.669676E-5   -3.255764E-6   3.255764E-6   -5.669676E-5   5.679017E-5   -1.767134E+2   -8.671345E+1   
4.470644E+3   8.003790E+1   8.003790E+1   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.150000E+3   -1.150000E+3   -4.060909E-2   5.091013E-2   -5.826367E-5   -3.247860E-6   3.247860E-6   -5.826367E-5   5.835412E-5   -1.768094E+2   -8.680940E+1   
4.492717E+3   8.004379E+1   8.004379E+1   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.100000E+3   -1.100000E+3   -4.189024E-2   5.112179E-2   -5.919359E-5   -2.438662E-6   2.438662E-6   -5.919359E-5   5.924380E-5   -1.776409E+2   -8.764086E+1   
4.514791E+3   8.002859E+1   8.002859E+1   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   -4.348928E-2   5.361236E-2   -6.180426E-5   -2.884224E-6   2.884224E-6   -6.180426E-5   6.187153E-5   -1.773281E+2   -8.732811E+1   
4.536842E+3   8.003060E+1   8.003060E+1   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   -4.408201E-2   5.566420E-2   -6.350707E-5   -3.787256E-6   3.787256E-6   -6.350707E-5   6.361989E-5   -1.765872E+2   -8.658720E+1   
4.558773E+3   7.995880E+1   7.995880E+1   -9.500000E+2   -9.500000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   -4.572276E-2   5.758533E-2   -6.577266E-5   -3.829691E-6   3.829691E-6   -6.577266E-5   6.588406E-5   -1.766676E+2   -8.666765E+1   
4.580443E+3   8.003301E+1   8.003301E+1   -9.000000E+2   -9.000000E+2   9.000000E+1   -8.990000E+2   -8.990000E+2   -4.686651E-2   5.948132E-2   -6.771462E-5   -4.223281E-6   4.223281E-6   -6.771462E-5   6.784619E-5   -1.764312E+2   -8.643115E+1   
4.602371E+3   7.997390E+1   7.997390E+1   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   -4.885334E-2   6.052195E-2   -6.962072E-5   -3.434091E-6   3.434091E-6   -6.962072E-5   6.970537E-5   -1.771761E+2   -8.717613E+1   
4.624095E+3   8.003188E+1   8.003188E+1   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   -4.911290E-2   6.280510E-2   -7.126819E-5   -4.734773E-6   4.734773E-6   -7.126819E-5   7.142530E-5   -1.761991E+2   -8.619908E+1   
4.645804E+3   8.006451E+1   8.006451E+1   -7.510000E+2   -7.510000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   -5.028241E-2   6.482686E-2   -7.330798E-5   -5.191541E-6   5.191541E-6   -7.330798E-5   7.349158E-5   -1.759492E+2   -8.594918E+1   
4.667786E+3   8.004559E+1   8.004559E+1   -7.000000E+2   -7.000000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   -5.065611E-2   6.532264E-2   -7.386192E-5   -5.239266E-6   5.239266E-6   -7.386192E-5   7.404750E-5   -1.759426E+2   -8.594262E+1   
4.689625E+3   8.000939E+1   8.000939E+1   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.490000E+2   -6.490000E+2   -5.289873E-2   6.870470E-2   -7.745111E-5   -5.791643E-6   5.791643E-6   -7.745111E-5   7.766736E-5   -1.757235E+2   -8.572349E+1   
4.711239E+3   8.004330E+1   8.004330E+1   -6.000000E+2   -6.000000E+2   9.000000E+1   -6.000000E+2   -6.000000E+2   -5.299816E-2   6.976621E-2   -7.820394E-5   -6.412096E-6   6.412096E-6   -7.820394E-5   7.846637E-5   -1.753127E+2   -8.531269E+1   
4.732976E+3   8.002841E+1   8.002841E+1   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   -5.524205E-2   7.092958E-2   -8.034890E-5   -5.513021E-6   5.513021E-6   -8.034890E-5   8.053781E-5   -1.760749E+2   -8.607489E+1   
4.754640E+3   8.000579E+1   8.000579E+1   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   -5.614400E-2   7.279610E-2   -8.212217E-5   -6.066188E-6   6.066188E-6   -8.212217E-5   8.234592E-5   -1.757754E+2   -8.577536E+1   
4.776368E+3   8.005441E+1   8.005441E+1   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   -5.698461E-2   7.432454E-2   -8.363734E-5   -6.443698E-6   6.443698E-6   -8.363734E-5   8.388520E-5   -1.755944E+2   -8.559445E+1   
4.797994E+3   8.000891E+1   8.000891E+1   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   -5.936534E-2   7.570450E-2   -8.600796E-5   -5.585016E-6   5.585016E-6   -8.600796E-5   8.618911E-5   -1.762847E+2   -8.628466E+1   
4.819690E+3   8.000259E+1   8.000259E+1   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   -5.985866E-2   7.816803E-2   -8.791743E-5   -6.830730E-6   6.830730E-6   -8.791743E-5   8.818239E-5   -1.755573E+2   -8.555734E+1   
4.841302E+3   8.002291E+1   8.002291E+1   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   -6.064710E-2   7.971916E-2   -8.941512E-5   -7.261661E-6   7.261661E-6   -8.941512E-5   8.970950E-5   -1.753570E+2   -8.535703E+1   
4.862939E+3   8.000820E+1   8.000820E+1   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   -6.222588E-2   8.043585E-2   -9.085797E-5   -6.562499E-6   6.562499E-6   -9.085797E-5   9.109466E-5   -1.758688E+2   -8.586881E+1   
4.884617E+3   8.001779E+1   8.001779E+1   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   -6.304623E-2   8.217108E-2   -9.249528E-5   -7.090182E-6   7.090182E-6   -9.249528E-5   9.276663E-5   -1.756166E+2   -8.561659E+1   
4.906243E+3   8.003149E+1   8.003149E+1   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   -6.365490E-2   8.473524E-2   -9.454160E-5   -8.316361E-6   8.316361E-6   -9.454160E-5   9.490667E-5   -1.749729E+2   -8.497291E+1   
4.927837E+3   8.001110E+1   8.001110E+1   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   -6.567607E-2   8.619127E-2   -9.673948E-5   -7.773362E-6   7.773362E-6   -9.673948E-5   9.705129E-5   -1.754060E+2   -8.540595E+1   
4.949469E+3   8.005279E+1   8.005279E+1   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   -6.529134E-2   8.858548E-2   -9.806095E-5   -9.623183E-6   9.623183E-6   -9.806095E-5   9.853200E-5   -1.743952E+2   -8.439524E+1   
4.982515E+3   7.999539E+1   7.999539E+1   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.600000E+1   -4.600000E+1   -6.687315E-2   8.835970E-2   -9.889185E-5   -8.305620E-6   8.305620E-6   -9.889185E-5   9.924002E-5   -1.751992E+2   -8.519917E+1   
5.004808E+3   8.004150E+1   8.004150E+1   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   -6.653692E-2   8.798049E-2   -9.843700E-5   -8.306392E-6   8.306392E-6   -9.843700E-5   9.878683E-5   -1.751766E+2   -8.517665E+1   
5.027035E+3   8.002700E+1   8.002700E+1   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   -6.682959E-2   8.804308E-2   -9.865871E-5   -8.130839E-6   8.130839E-6   -9.865871E-5   9.899319E-5   -1.752887E+2   -8.528868E+1   
5.049227E+3   8.000131E+1   8.000131E+1   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   -6.650439E-2   8.881558E-2   -9.896077E-5   -8.876408E-6   8.876408E-6   -9.896077E-5   9.935807E-5   -1.748745E+2   -8.487450E+1   
5.071463E+3   8.004391E+1   8.004391E+1   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   -6.700569E-2   8.768228E-2   -9.853259E-5   -7.764710E-6   7.764710E-6   -9.853259E-5   9.883806E-5   -1.754942E+2   -8.549421E+1   
5.093734E+3   8.005230E+1   8.005230E+1   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   -6.719959E-2   8.775225E-2   -9.869803E-5   -7.667038E-6   7.667038E-6   -9.869803E-5   9.899538E-5   -1.755581E+2   -8.555808E+1   
5.115989E+3   8.000439E+1   8.000439E+1   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   -6.654367E-2   8.899353E-2   -9.910095E-5   -8.963692E-6   8.963692E-6   -9.910095E-5   9.950551E-5   -1.748317E+2   -8.483165E+1   
5.138279E+3   7.999828E+1   7.999828E+1   -3.300000E+1   -3.300000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   -6.775242E-2   8.786758E-2   -9.911494E-5   -7.333546E-6   7.333546E-6   -9.911494E-5   9.938588E-5   -1.757684E+2   -8.576838E+1   
5.159519E+3   8.002691E+1   8.002691E+1   -3.100000E+1   -3.100000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   -6.683389E-2   8.829649E-2   -9.882641E-5   -8.293329E-6   8.293329E-6   -9.882641E-5   9.917378E-5   -1.752031E+2   -8.520308E+1   
5.180789E+3   8.000790E+1   8.000790E+1   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   -6.554414E-2   8.873703E-2   -9.831594E-5   -9.535288E-6   9.535288E-6   -9.831594E-5   9.877725E-5   -1.744604E+2   -8.446043E+1   
5.203073E+3   8.005950E+1   8.005950E+1   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.600000E+1   -2.600000E+1   -6.779291E-2   8.945494E-2   -1.001738E-4   -8.341367E-6   8.341367E-6   -1.001738E-4   1.005205E-4   -1.752400E+2   -8.524002E+1   
5.225298E+3   7.999630E+1   7.999630E+1   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   -6.750392E-2   8.920030E-2   -9.982929E-5   -8.388637E-6   8.388637E-6   -9.982929E-5   1.001811E-4   -1.751967E+2   -8.519673E+1   
5.247550E+3   8.003051E+1   8.003051E+1   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   -6.708853E-2   8.916840E-2   -9.955170E-5   -8.675019E-6   8.675019E-6   -9.955170E-5   9.992896E-5   -1.750198E+2   -8.501978E+1   
5.269810E+3   7.997231E+1   7.997231E+1   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   -6.779293E-2   8.826090E-2   -9.939614E-5   -7.560727E-6   7.560727E-6   -9.939614E-5   9.968329E-5   -1.756501E+2   -8.565008E+1   
5.292064E+3   7.998669E+1   7.998669E+1   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   -6.671976E-2   8.985131E-2   -9.976848E-5   -9.394245E-6   9.394245E-6   -9.976848E-5   1.002098E-4   -1.746209E+2   -8.462086E+1   
5.314333E+3   8.001730E+1   8.001730E+1   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   -6.793773E-2   8.962185E-2   -1.003720E-4   -8.343377E-6   8.343377E-6   -1.003720E-4   1.007182E-4   -1.752482E+2   -8.524824E+1   
5.336570E+3   8.001599E+1   8.001599E+1   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   -6.595645E-2   8.894014E-2   -9.870313E-5   -9.363110E-6   9.363110E-6   -9.870313E-5   9.914624E-5   -1.745811E+2   -8.458106E+1   
5.358861E+3   8.002041E+1   8.002041E+1   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   -6.753705E-2   8.953839E-2   -1.000700E-4   -8.585172E-6   8.585172E-6   -1.000700E-4   1.004376E-4   -1.750965E+2   -8.509650E+1   
5.381092E+3   8.000479E+1   8.000479E+1   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   -6.771867E-2   8.963103E-2   -1.002426E-4   -8.511404E-6   8.511404E-6   -1.002426E-4   1.006033E-4   -1.751468E+2   -8.514677E+1   
5.403279E+3   8.004449E+1   8.004449E+1   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   -6.796044E-2   8.951753E-2   -1.003181E-4   -8.258377E-6   8.258377E-6   -1.003181E-4   1.006575E-4   -1.752939E+2   -8.529392E+1   
5.425355E+3   8.002810E+1   8.002810E+1   -7.000000E+0   -7.000000E+0   9.000000E+1   -6.000000E+0   -6.000000E+0   -6.775918E-2   8.992802E-2   -1.004611E-4   -8.675608E-6   8.675608E-6   -1.004611E-4   1.008350E-4   -1.750643E+2   -8.506430E+1   
5.446442E+3   8.004989E+1   8.004989E+1   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   -6.807823E-2   8.951569E-2   -1.003898E-4   -8.170059E-6   8.170059E-6   -1.003898E-4   1.007217E-4   -1.753473E+2   -8.534733E+1   
5.468520E+3   8.006011E+1   8.006011E+1   -4.000000E+0   -4.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   -6.675044E-2   8.941260E-2   -9.950173E-5   -9.084734E-6   9.084734E-6   -9.950173E-5   9.991560E-5   -1.747832E+2   -8.478323E+1   
5.490527E+3   8.002361E+1   8.002361E+1   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   -6.678235E-2   8.921503E-2   -9.939278E-5   -8.931961E-6   8.931961E-6   -9.939278E-5   9.979331E-5   -1.748649E+2   -8.486489E+1   
5.512476E+3   8.002371E+1   8.002371E+1   0.000000E+0   0.000000E+0   9.000000E+1   0.000000E+0   0.000000E+0   -6.812731E-2   8.881495E-2   -9.996373E-5   -7.675634E-6   7.675634E-6   -9.996373E-5   1.002580E-4   -1.756092E+2   -8.560921E+1   
5.534460E+3   7.999200E+1   7.999200E+1   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   -6.861941E-2   8.873703E-2   -1.002172E-4   -7.260716E-6   7.260716E-6   -1.002172E-4   1.004799E-4   -1.758562E+2   -8.585617E+1   
5.555988E+3   7.999420E+1   7.999420E+1   3.000000E+0   3.000000E+0   9.000000E+1   3.000000E+0   3.000000E+0   -6.886731E-2   8.854315E-2   -1.002442E-4   -6.950611E-6   6.950611E-6   -1.002442E-4   1.004849E-4   -1.760336E+2   -8.603364E+1   
5.577676E+3   7.998950E+1   7.998950E+1   5.000000E+0   5.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   -6.869061E-2   9.008816E-2   -1.011412E-4   -8.091390E-6   8.091390E-6   -1.011412E-4   1.014644E-4   -1.754260E+2   -8.542603E+1   
5.599400E+3   8.003719E+1   8.003719E+1   7.000000E+0   7.000000E+0   9.000000E+1   7.000000E+0   7.000000E+0   -6.873048E-2   9.012745E-2   -1.011915E-4   -8.087587E-6   8.087587E-6   -1.011915E-4   1.015141E-4   -1.754304E+2   -8.543043E+1   
5.621130E+3   8.001519E+1   8.001519E+1   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   -6.912685E-2   8.916717E-2   -1.008111E-4   -7.166611E-6   7.166611E-6   -1.008111E-4   1.010655E-4   -1.759337E+2   -8.593371E+1   
5.643000E+3   8.002599E+1   8.002599E+1   1.100000E+1   1.100000E+1   9.000000E+1   1.100000E+1   1.100000E+1   -6.825434E-2   9.027163E-2   -1.009910E-4   -8.534007E-6   8.534007E-6   -1.009910E-4   1.013509E-4   -1.751698E+2   -8.516983E+1   
5.665078E+3   8.000649E+1   8.000649E+1   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   -6.786041E-2   9.003662E-2   -1.005944E-4   -8.671729E-6   8.671729E-6   -1.005944E-4   1.009675E-4   -1.750730E+2   -8.507300E+1   
5.686979E+3   8.004241E+1   8.004241E+1   1.500000E+1   1.500000E+1   9.000000E+1   1.500000E+1   1.500000E+1   -6.885566E-2   8.867201E-2   -1.003209E-4   -7.043474E-6   7.043474E-6   -1.003209E-4   1.005679E-4   -1.759839E+2   -8.598389E+1   
5.708992E+3   8.001150E+1   8.001150E+1   1.700000E+1   1.700000E+1   9.000000E+1   1.700000E+1   1.700000E+1   -6.855560E-2   8.985194E-2   -1.009039E-4   -8.036804E-6   8.036804E-6   -1.009039E-4   1.012234E-4   -1.754461E+2   -8.544611E+1   
5.731007E+3   7.999789E+1   7.999789E+1   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   -6.791136E-2   9.010349E-2   -1.006694E-4   -8.677766E-6   8.677766E-6   -1.006694E-4   1.010427E-4   -1.750732E+2   -8.507325E+1   
5.752843E+3   7.998589E+1   7.998589E+1   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   -6.835126E-2   8.995562E-2   -1.008451E-4   -8.255728E-6   8.255728E-6   -1.008451E-4   1.011825E-4   -1.753199E+2   -8.531989E+1   
5.774710E+3   8.003661E+1   8.003661E+1   2.300000E+1   2.300000E+1   9.000000E+1   2.300000E+1   2.300000E+1   -6.895628E-2   9.098893E-2   -1.018921E-4   -8.483781E-6   8.483781E-6   -1.018921E-4   1.022447E-4   -1.752404E+2   -8.524040E+1   
5.796837E+3   7.998489E+1   7.998489E+1   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   -6.702655E-2   9.099690E-2   -1.007043E-4   -9.916282E-6   9.916282E-6   -1.007043E-4   1.011913E-4   -1.743763E+2   -8.437625E+1   
5.818782E+3   7.997411E+1   7.997411E+1   2.600000E+1   2.600000E+1   9.000000E+1   2.700000E+1   2.700000E+1   -6.894156E-2   9.091716E-2   -1.018363E-4   -8.447751E-6   8.447751E-6   -1.018363E-4   1.021861E-4   -1.752579E+2   -8.525793E+1   
5.840661E+3   8.006530E+1   8.006530E+1   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   -6.933855E-2   9.033300E-2   -1.017013E-4   -7.772218E-6   7.772218E-6   -1.017013E-4   1.019978E-4   -1.756298E+2   -8.562983E+1   
5.862542E+3   8.000079E+1   8.000079E+1   3.100000E+1   3.100000E+1   9.000000E+1   3.100000E+1   3.100000E+1   -6.965148E-2   9.117236E-2   -1.024414E-4   -8.089515E-6   8.089515E-6   -1.024414E-4   1.027603E-4   -1.754849E+2   -8.548488E+1   
5.884679E+3   8.001599E+1   8.001599E+1   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   -6.761684E-2   9.190871E-2   -1.016631E-4   -1.007580E-5   1.007580E-5   -1.016631E-4   1.021611E-4   -1.743399E+2   -8.433991E+1   
5.906615E+3   8.002679E+1   8.002679E+1   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   -6.856910E-2   9.074837E-2   -1.014961E-4   -8.612884E-6   8.612884E-6   -1.014961E-4   1.018609E-4   -1.751495E+2   -8.514954E+1   
5.928553E+3   8.001879E+1   8.001879E+1   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   -7.021105E-2   9.139452E-2   -1.029320E-4   -7.820876E-6   7.820876E-6   -1.029320E-4   1.032287E-4   -1.756550E+2   -8.565496E+1   
5.950445E+3   8.000939E+1   8.000939E+1   3.900000E+1   3.900000E+1   9.000000E+1   3.900000E+1   3.900000E+1   -6.822428E-2   9.121473E-2   -1.015866E-4   -9.172820E-6   9.172820E-6   -1.015866E-4   1.019999E-4   -1.748404E+2   -8.484044E+1   
5.972503E+3   8.003631E+1   8.003631E+1   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   -6.899554E-2   9.151354E-2   -1.022581E-4   -8.797729E-6   8.797729E-6   -1.022581E-4   1.026358E-4   -1.750827E+2   -8.508269E+1   
5.994345E+3   8.002831E+1   8.002831E+1   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   -6.924958E-2   9.132520E-2   -1.022925E-4   -8.486695E-6   8.486695E-6   -1.022925E-4   1.026439E-4   -1.752573E+2   -8.525732E+1   
6.016276E+3   8.001730E+1   8.001730E+1   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   -6.944777E-2   9.073121E-2   -1.020281E-4   -7.951772E-6   7.951772E-6   -1.020281E-4   1.023375E-4   -1.755435E+2   -8.554354E+1   
6.038211E+3   8.001971E+1   8.001971E+1   4.700000E+1   4.700000E+1   9.000000E+1   4.800000E+1   4.800000E+1   -6.883173E-2   9.073367E-2   -1.016489E-4   -8.409026E-6   8.409026E-6   -1.016489E-4   1.019961E-4   -1.752709E+2   -8.527091E+1   
6.060332E+3   8.002450E+1   8.002450E+1   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   -6.911460E-2   9.081715E-2   -1.018781E-4   -8.254386E-6   8.254386E-6   -1.018781E-4   1.022120E-4   -1.753679E+2   -8.536789E+1   
6.094200E+3   8.004501E+1   8.004501E+1   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   -7.157322E-2   9.289969E-2   -1.047545E-4   -7.797419E-6   7.797419E-6   -1.047545E-4   1.050443E-4   -1.757430E+2   -8.574303E+1   
6.116544E+3   8.000799E+1   8.000799E+1   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   -7.153517E-2   9.590276E-2   -1.066868E-4   -9.788881E-6   9.788881E-6   -1.066868E-4   1.071350E-4   -1.747576E+2   -8.475760E+1   
6.138928E+3   8.006170E+1   8.006170E+1   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   -7.190333E-2   9.650842E-2   -1.073089E-4   -9.912542E-6   9.912542E-6   -1.073089E-4   1.077658E-4   -1.747223E+2   -8.472234E+1   
6.161305E+3   7.999740E+1   7.999740E+1   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   -7.376127E-2   9.783685E-2   -1.093228E-4   -9.406840E-6   9.406840E-6   -1.093228E-4   1.097267E-4   -1.750820E+2   -8.508201E+1   
6.183936E+3   8.001949E+1   8.001949E+1   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   -7.575418E-2   9.912417E-2   -1.113933E-4   -8.774437E-6   8.774437E-6   -1.113933E-4   1.117383E-4   -1.754961E+2   -8.549612E+1   
6.206276E+3   8.002239E+1   8.002239E+1   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   -7.727220E-2   1.004925E-1   -1.132230E-4   -8.546210E-6   8.546210E-6   -1.132230E-4   1.135450E-4   -1.756834E+2   -8.568343E+1   
6.228592E+3   8.000469E+1   8.000469E+1   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   -7.762133E-2   1.029621E-1   -1.150473E-4   -9.902590E-6   9.902590E-6   -1.150473E-4   1.154727E-4   -1.750804E+2   -8.508044E+1   
6.251476E+3   8.000591E+1   8.000591E+1   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   -7.970630E-2   1.038193E-1   -1.168946E-4   -8.920886E-6   8.920886E-6   -1.168946E-4   1.172345E-4   -1.756359E+2   -8.563589E+1   
6.273704E+3   7.998510E+1   7.998510E+1   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   -7.967990E-2   1.073554E-1   -1.191813E-4   -1.125220E-5   1.125220E-5   -1.191813E-4   1.197113E-4   -1.746066E+2   -8.460655E+1   
6.296341E+3   8.000869E+1   8.000869E+1   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   -8.068066E-2   1.078812E-1   -1.201425E-4   -1.085578E-5   1.085578E-5   -1.201425E-4   1.206319E-4   -1.748369E+2   -8.483691E+1   
6.319628E+3   8.001440E+1   8.001440E+1   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   -8.368354E-2   1.096349E-1   -1.231411E-4   -9.781233E-6   9.781233E-6   -1.231411E-4   1.235290E-4   -1.754585E+2   -8.545847E+1   
6.342235E+3   8.003051E+1   8.003051E+1   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   -8.444440E-2   1.116118E-1   -1.248991E-4   -1.051096E-5   1.051096E-5   -1.248991E-4   1.253406E-4   -1.751896E+2   -8.518957E+1   
6.364865E+3   8.003610E+1   8.003610E+1   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   -8.437567E-2   1.131446E-1   -1.258549E-4   -1.156386E-5   1.156386E-5   -1.258549E-4   1.263850E-4   -1.747503E+2   -8.475026E+1   
6.388280E+3   8.001150E+1   8.001150E+1   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   -8.754239E-2   1.143896E-1   -1.286235E-4   -1.003560E-5   1.003560E-5   -1.286235E-4   1.290144E-4   -1.755386E+2   -8.553865E+1   
6.410854E+3   8.001690E+1   8.001690E+1   7.980000E+2   7.980000E+2   9.000000E+1   7.980000E+2   7.980000E+2   -8.793388E-2   1.167359E-1   -1.303937E-4   -1.128001E-5   1.128001E-5   -1.303937E-4   1.308807E-4   -1.750558E+2   -8.505580E+1   
6.433442E+3   8.003369E+1   8.003369E+1   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   -8.956417E-2   1.182564E-1   -1.323919E-4   -1.106823E-5   1.106823E-5   -1.323919E-4   1.328537E-4   -1.752211E+2   -8.522107E+1   
6.456741E+3   8.003741E+1   8.003741E+1   8.980000E+2   8.980000E+2   9.000000E+1   8.980000E+2   8.980000E+2   -9.359004E-2   1.219416E-1   -1.372810E-4   -1.049985E-5   1.049985E-5   -1.372810E-4   1.376819E-4   -1.756263E+2   -8.562629E+1   
6.479342E+3   8.001190E+1   8.001190E+1   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   -9.637029E-2   1.253371E-1   -1.412114E-4   -1.066342E-5   1.066342E-5   -1.412114E-4   1.416134E-4   -1.756816E+2   -8.568157E+1   
6.501924E+3   8.004470E+1   8.004470E+1   9.980000E+2   9.980000E+2   9.000000E+1   9.980000E+2   9.980000E+2   -9.771716E-2   1.279510E-1   -1.437465E-4   -1.137611E-5   1.137611E-5   -1.437465E-4   1.441959E-4   -1.754750E+2   -8.547504E+1   
6.525455E+3   8.002981E+1   8.002981E+1   1.047000E+3   1.047000E+3   9.000000E+1   1.048000E+3   1.048000E+3   -9.987335E-2   1.283425E-1   -1.453345E-4   -1.003726E-5   1.003726E-5   -1.453345E-4   1.456807E-4   -1.760492E+2   -8.604924E+1   
6.548259E+3   8.002001E+1   8.002001E+1   1.098000E+3   1.098000E+3   9.000000E+1   1.098000E+3   1.098000E+3   -9.776011E-2   1.306189E-1   -1.455106E-4   -1.308851E-5   1.308851E-5   -1.455106E-4   1.460980E-4   -1.748601E+2   -8.486014E+1   
6.571146E+3   8.003781E+1   8.003781E+1   1.148000E+3   1.148000E+3   9.000000E+1   1.148000E+3   1.148000E+3   -1.010809E-1   1.314325E-1   -1.480935E-4   -1.116428E-5   1.116428E-5   -1.480935E-4   1.485137E-4   -1.756888E+2   -8.568881E+1   
6.594637E+3   8.003851E+1   8.003851E+1   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   -1.017785E-1   1.330959E-1   -1.496082E-4   -1.173578E-5   1.173578E-5   -1.496082E-4   1.500678E-4   -1.755147E+2   -8.551471E+1   
6.617529E+3   7.997631E+1   7.997631E+1   1.248000E+3   1.248000E+3   9.000000E+1   1.248000E+3   1.248000E+3   -1.031223E-1   1.351079E-1   -1.517494E-4   -1.205726E-5   1.205726E-5   -1.517494E-4   1.522276E-4   -1.754571E+2   -8.545710E+1   
6.640317E+3   8.004312E+1   8.004312E+1   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   -1.035328E-1   1.367928E-1   -1.531005E-4   -1.285519E-5   1.285519E-5   -1.531005E-4   1.536392E-4   -1.752004E+2   -8.520038E+1   
6.663589E+3   8.002471E+1   8.002471E+1   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   -1.045771E-1   1.387826E-1   -1.550421E-4   -1.338370E-5   1.338370E-5   -1.550421E-4   1.556187E-4   -1.750663E+2   -8.506629E+1   
6.686163E+3   8.006341E+1   8.006341E+1   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   -1.070726E-1   1.401693E-1   -1.574881E-4   -1.244455E-5   1.244455E-5   -1.574881E-4   1.579790E-4   -1.754819E+2   -8.548193E+1   
6.708727E+3   8.001110E+1   8.001110E+1   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   -1.086255E-1   1.408872E-1   -1.589157E-4   -1.176527E-5   1.176527E-5   -1.589157E-4   1.593507E-4   -1.757659E+2   -8.576585E+1   
6.731758E+3   7.999749E+1   7.999749E+1   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   -1.094600E-1   1.441098E-1   -1.615305E-4   -1.325488E-5   1.325488E-5   -1.615305E-4   1.620734E-4   -1.753089E+2   -8.530893E+1   
6.754335E+3   7.998721E+1   7.998721E+1   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   -1.121942E-1   1.459524E-1   -1.644209E-4   -1.243725E-5   1.243725E-5   -1.644209E-4   1.648906E-4   -1.756742E+2   -8.567423E+1   
6.776865E+3   8.003570E+1   8.003570E+1   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   -1.117806E-1   1.484803E-1   -1.658117E-4   -1.439585E-5   1.439585E-5   -1.658117E-4   1.664354E-4   -1.750380E+2   -8.503799E+1   
6.799656E+3   8.005691E+1   8.005691E+1   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   -1.141177E-1   1.494228E-1   -1.678704E-4   -1.328338E-5   1.328338E-5   -1.678704E-4   1.683951E-4   -1.754757E+2   -8.547568E+1   
6.822186E+3   8.001821E+1   8.001821E+1   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   -1.153817E-1   1.522177E-1   -1.704721E-4   -1.417572E-5   1.417572E-5   -1.704721E-4   1.710605E-4   -1.752465E+2   -8.524647E+1   
6.844719E+3   8.000579E+1   8.000579E+1   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   -1.168261E-1   1.529190E-1   -1.718219E-4   -1.356591E-5   1.356591E-5   -1.718219E-4   1.723566E-4   -1.754857E+2   -8.548567E+1   
6.867539E+3   8.007610E+1   8.007610E+1   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   -1.176649E-1   1.536105E-1   -1.727908E-4   -1.339762E-5   1.339762E-5   -1.727908E-4   1.733094E-4   -1.755663E+2   -8.556635E+1   
6.890147E+3   7.999941E+1   7.999941E+1   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   -1.190976E-1   1.560784E-1   -1.752839E-4   -1.395134E-5   1.395134E-5   -1.752839E-4   1.758382E-4   -1.754493E+2   -8.544926E+1   
6.912658E+3   8.001269E+1   8.001269E+1   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   -1.219072E-1   1.589389E-1   -1.788840E-4   -1.374341E-5   1.374341E-5   -1.788840E-4   1.794111E-4   -1.756067E+2   -8.560667E+1   
6.935442E+3   8.001400E+1   8.001400E+1   1.949000E+3   1.949000E+3   9.000000E+1   1.949000E+3   1.949000E+3   -1.215059E-1   1.591837E-1   -1.787953E-4   -1.420027E-5   1.420027E-5   -1.787953E-4   1.793583E-4   -1.754590E+2   -8.545899E+1   
6.957973E+3   8.007241E+1   8.007241E+1   1.999000E+3   1.999000E+3   9.000000E+1   2.000000E+3   2.000000E+3   -1.208942E-1   1.612098E-1   -1.797366E-4   -1.597733E-5   1.597733E-5   -1.797366E-4   1.804454E-4   -1.749202E+2   -8.492016E+1   
6.995911E+3   8.004510E+1   8.004510E+1   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   -1.355766E-1   1.794596E-1   -2.007000E-4   -1.704895E-5   1.704895E-5   -2.007000E-4   2.014228E-4   -1.751445E+2   -8.514453E+1   
7.022524E+3   8.002111E+1   8.002111E+1   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   -1.509157E-1   1.990270E-1   -2.229273E-4   -1.849632E-5   1.849632E-5   -2.229273E-4   2.236933E-4   -1.752570E+2   -8.525702E+1   
7.048215E+3   8.004531E+1   8.004531E+1   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -1.681942E-1   2.227764E-1   -2.490774E-4   -2.124326E-5   2.124326E-5   -2.490774E-4   2.499817E-4   -1.751252E+2   -8.512517E+1   
7.074055E+3   8.000970E+1   8.000970E+1   3.999000E+3   3.999000E+3   9.000000E+1   4.000000E+3   4.000000E+3   -1.769519E-1   2.368895E-1   -2.636835E-4   -2.399252E-5   2.399252E-5   -2.636835E-4   2.647728E-4   -1.748010E+2   -8.480098E+1   
7.100699E+3   8.001531E+1   8.001531E+1   4.498000E+3   4.498000E+3   9.000000E+1   4.499000E+3   4.499000E+3   -1.878348E-1   2.526046E-1   -2.806470E-4   -2.621735E-5   2.621735E-5   -2.806470E-4   2.818689E-4   -1.746631E+2   -8.466306E+1   
7.126628E+3   8.003039E+1   8.003039E+1   4.998000E+3   4.998000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -1.953700E-1   2.637553E-1   -2.925679E-4   -2.793402E-5   2.793402E-5   -2.925679E-4   2.938984E-4   -1.745460E+2   -8.454600E+1   
7.152381E+3   8.001891E+1   8.001891E+1   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -1.939293E-1   2.640075E-1   -2.918415E-4   -2.916454E-5   2.916454E-5   -2.918415E-4   2.932951E-4   -1.742932E+2   -8.429322E+1   
7.178783E+3   8.006509E+1   8.006509E+1   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -1.792296E-1   2.495355E-1   -2.733279E-4   -3.057547E-5   3.057547E-5   -2.733279E-4   2.750327E-4   -1.736172E+2   -8.361722E+1   
7.204727E+3   8.003289E+1   8.003289E+1   6.498000E+3   6.498000E+3   9.000000E+1   6.499000E+3   6.499000E+3   -1.685133E-1   2.354389E-1   -2.575217E-4   -2.928568E-5   2.928568E-5   -2.575217E-4   2.591815E-4   -1.735121E+2   -8.351213E+1   
7.230877E+3   8.002401E+1   8.002401E+1   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -1.574448E-1   2.240809E-1   -2.432813E-4   -3.004666E-5   3.004666E-5   -2.432813E-4   2.451297E-4   -1.729593E+2   -8.295929E+1   
7.256559E+3   7.999490E+1   7.999490E+1   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -1.519925E-1   2.189906E-1   -2.365951E-4   -3.075147E-5   3.075147E-5   -2.365951E-4   2.385852E-4   -1.725945E+2   -8.259449E+1   
7.282044E+3   8.001199E+1   8.001199E+1   7.999000E+3   7.999000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -1.503180E-1   2.202227E-1   -2.363623E-4   -3.279546E-5   3.279546E-5   -2.363623E-4   2.386267E-4   -1.721006E+2   -8.210060E+1   
7.308436E+3   8.005721E+1   8.005721E+1   8.498000E+3   8.498000E+3   9.000000E+1   8.499000E+3   8.499000E+3   -1.507666E-1   2.272451E-1   -2.412133E-4   -3.705481E-5   3.705481E-5   -2.412133E-4   2.440428E-4   -1.712666E+2   -8.126658E+1   
7.334878E+3   8.000741E+1   8.000741E+1   8.998000E+3   8.998000E+3   9.000000E+1   8.999000E+3   8.999000E+3   -1.681967E-1   2.458012E-1   -2.640748E-4   -3.629440E-5   3.629440E-5   -2.640748E-4   2.665573E-4   -1.721743E+2   -8.217431E+1   
7.361264E+3   7.999090E+1   7.999090E+1   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -1.798542E-1   2.615250E-1   -2.815227E-4   -3.795185E-5   3.795185E-5   -2.815227E-4   2.840693E-4   -1.723223E+2   -8.232229E+1   
7.386641E+3   8.003561E+1   8.003561E+1   9.998000E+3   9.998000E+3   9.000000E+1   1.000000E+4   1.000000E+4   -1.888872E-1   2.786157E-1   -2.982384E-4   -4.244428E-5   4.244428E-5   -2.982384E-4   3.012435E-4   -1.719002E+2   -8.190025E+1   
@@END Data.
@Time at end of measurement: 12:52:32
@NO Instrument  Changes.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -9499.000      -9999.000      250.000        Coercive Field: Field at which M//H changes sign
Ms  emu                                 3.260E-4       -3.982E-4      3.621E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -9.996E-5      1.375E-4       1.187E-4       Remanent Magnetization: M at H=0        
S                                       0.307          0.345          0.326          Squareness: Mr/Ms                       
S*                                      1.223          1.245          1.234          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
