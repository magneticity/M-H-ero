@Filename: c:\vsm-lv\Will\data\AJA335e-FePtFeRh_1030nm_Tann_6\AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_100deg.VHD
@Measurement Controlfilename: C:\vsm-lv\Will\Recipes\10kOe OoP loop 100deg.VHC
@Signal Manipulation filename: c:\vsm-lv\Will\settings\default.cal
@Operator: Will
@Samplename: AJA335e-FePtFeRh_1030nm_Tann_6
@Date: 07 November 2019    (2019-07-11)
@Time: 15:14:47
@Test ID: AJA335e-FePtFeRh_1030nm_Tann_600deg_OoP_100deg
@Apparatus: DMS Model 10; SN:20090630; Customer: Manchester; first started on: Monday, August 24, 2009
VSM Model = DMS Model 10, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 10 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = DMS Rotating Base
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = E-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = TRUE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = TRUE, Sensor Angle = 45 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: DMS EasyVSM Software version 9.12f (June 2, 2009)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 90.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 1:      Set Sample Temperature to 100.1270 [degC] and wait 60.0000 s ; Set Mode = Set and wait till there
Action 2:      Set Applied Field to 9999.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there
Action 3:      Set Auto Range Signal to 13.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 5
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 5.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: 10000.0000 [Oe] To: 2000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Measured Signal(s) = Parallel & Perpendicular to Sample
@Section 0 END
@Section 1: Hysteresis
@Main Parameter Setup:
     From: 2000.0000 [Oe] To: 50.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: 50.0000 [Oe] To: -50.0000 [Oe] Min Stepsize/Sweeprate =  2.0000 [Oe] Max Stepsize/Sweeprate =  2.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Main Parameter Setup:
     From: -50.0000 [Oe] To: -2000.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Main Parameter Setup:
     From: -2000.0000 [Oe] To: -10000.0000 [Oe] Min Stepsize/Sweeprate = 500.0000 [Oe] Max Stepsize/Sweeprate = 500.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    5.00 [sec] Up & Down = No
@Section 4 END
@@Plot Settings
Number of plots: 2
Plot 0: Hysteresis = On; Section: 0; Signal: Parallel with Sample; Label: Hys Parallel with Sample; Point style: 2; Interpolation: On; Color: 0; Mirror: Off
Plot 1: Hysteresis = On; Section: 0; Signal: Perpendicular to Sample; Label: Hys Perp to Sample; Point style: 0; Interpolation: On; Color: 16740729; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = TRUE
Sensor Angle = 45 deg
@Gauss Range: 30 kOe
@Emu Range: 50 uV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 75
@Rot 0 deg cal: -21100
@Rot 360 deg cal: 20910
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 24.706
@Y Coils Correction Factor: 0.964
@Sample Shape Correction Factor: 0.919
@Coil Angle Alpha: 42.300
@Coil Angle Beta: -47.320
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
15000.000000   1.000000
15249.000000   1.000524
15499.000000   1.000702
15750.000000   1.001233
16000.000000   1.001406
16250.000000   1.001585
16499.000000   1.001758
16749.000000   1.001937
16999.000000   1.002110
17249.000000   1.001937
17499.000000   1.002289
17749.000000   1.002289
17999.000000   1.002289
18249.000000   1.002462
18499.000000   1.002462
18748.000000   1.002462
18999.000000   1.002462
19249.000000   1.002462
19499.000000   1.002642
19749.000000   1.002642
19999.000000   1.002462
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = No
Angular Sensitivity Correction = No
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = 25 October 2019  12:02:56
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 5
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Raw Applied Field, Applied Field [Oe]
Column 4: Applied Field, Applied Field [Oe]
Column 5: Field Angle, Field Angle [deg]
Column 6: Raw Applied Field For Plot , Applied Field [Oe]
Column 7: Applied Field For Plot , Applied Field [Oe]
Column 8: Raw Signal Mx, Moment as measured [memu]
Column 9: Raw Signal My, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
Column 11: Signal Y direction, Moment [emu]
Column 12: Signal parallel with sample, Moment [emu]
Column 13: Signal perpendicular to sample, Moment [emu]
Column 14: Signal Magnitude, Moment [emu]
Column 15: Signal Angle with field, Angle [deg]
Column 16: Signal Angle with sample, Angle [deg]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Raw_Signal_My   Signal_X_direction   Signal_Y_direction   Signal_parallel_with_sample   Signal_perpendicular_to_sample   Signal_Magnitude   Signal_Angle_with_field   Signal_Angle_with_sample      
@Time at start of measurement: 15:14:47
@@Data
New Section: Section 0: 
3.211600E+1   1.000335E+2   1.000335E+2   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -2.402697E-1   3.221747E-1   -3.583749E-4   -3.291777E-5   3.291777E-5   -3.583749E-4   3.598835E-4   -1.747519E+2   -8.475194E+1   
5.749200E+1   9.994659E+1   9.994659E+1   9.498000E+3   9.498000E+3   9.000000E+1   9.498000E+3   9.498000E+3   -2.210013E-1   2.970521E-1   -3.301002E-4   -3.074484E-5   3.074484E-5   -3.301002E-4   3.315289E-4   -1.746789E+2   -8.467894E+1   
8.255700E+1   1.000198E+2   1.000198E+2   8.998000E+3   8.998000E+3   9.000000E+1   8.998000E+3   8.998000E+3   -1.984085E-1   2.707434E-1   -2.989977E-4   -3.025533E-5   3.025533E-5   -2.989977E-4   3.005246E-4   -1.742220E+2   -8.422196E+1   
1.077000E+2   1.000381E+2   1.000381E+2   8.497000E+3   8.497000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -1.751695E-1   2.443390E-1   -2.674334E-4   -3.018118E-5   3.018118E-5   -2.674334E-4   2.691310E-4   -1.735611E+2   -8.356113E+1   
1.337120E+2   1.000746E+2   1.000746E+2   7.999000E+3   7.999000E+3   9.000000E+1   7.999000E+3   7.999000E+3   -1.547561E-1   2.189004E-1   -2.382450E-4   -2.864849E-5   2.864849E-5   -2.382450E-4   2.399612E-4   -1.731432E+2   -8.314322E+1   
1.595560E+2   1.000460E+2   1.000460E+2   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -1.330873E-1   1.928548E-1   -2.078851E-4   -2.764753E-5   2.764753E-5   -2.078851E-4   2.097155E-4   -1.724244E+2   -8.242444E+1   
1.851370E+2   1.000075E+2   1.000075E+2   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -1.113946E-1   1.672769E-1   -1.778151E-4   -2.696997E-5   2.696997E-5   -1.778151E-4   1.798488E-4   -1.713754E+2   -8.137544E+1   
2.105520E+2   9.999371E+1   9.999371E+1   6.497000E+3   6.497000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -9.545969E-2   1.465666E-1   -1.544749E-4   -2.521613E-5   2.521613E-5   -1.544749E-4   1.565195E-4   -1.707289E+2   -8.072894E+1   
2.360230E+2   1.000431E+2   1.000431E+2   5.998000E+3   5.998000E+3   9.000000E+1   5.998000E+3   5.998000E+3   -7.650768E-2   1.212304E-1   -1.262567E-4   -2.266957E-5   2.266957E-5   -1.262567E-4   1.282757E-4   -1.698209E+2   -7.982092E+1   
2.618590E+2   1.000793E+2   1.000793E+2   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -6.173683E-2   1.025498E-1   -1.049582E-4   -2.138169E-5   2.138169E-5   -1.049582E-4   1.071140E-4   -1.684855E+2   -7.848548E+1   
2.872160E+2   1.000172E+2   1.000172E+2   4.997000E+3   4.997000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -4.564912E-2   8.287486E-2   -8.219794E-5   -2.041774E-5   2.041774E-5   -8.219794E-5   8.469584E-5   -1.660502E+2   -7.605022E+1   
3.123510E+2   9.997979E+1   9.997979E+1   4.498000E+3   4.498000E+3   9.000000E+1   4.498000E+3   4.498000E+3   -2.867239E-2   5.954204E-2   -5.650571E-5   -1.771991E-5   1.771991E-5   -5.650571E-5   5.921901E-5   -1.625888E+2   -7.258883E+1   
3.382060E+2   1.000365E+2   1.000365E+2   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -1.727313E-2   4.083980E-2   -3.727758E-5   -1.392417E-5   1.392417E-5   -3.727758E-5   3.979322E-5   -1.595180E+2   -6.951801E+1   
3.635470E+2   1.000289E+2   1.000289E+2   3.498000E+3   3.498000E+3   9.000000E+1   3.498000E+3   3.498000E+3   6.356788E-4   2.015208E-2   -1.273183E-5   -1.364503E-5   1.364503E-5   -1.273183E-5   1.866243E-5   -1.330171E+2   -4.301714E+1   
3.889050E+2   1.000666E+2   1.000666E+2   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   1.510778E-2   3.067947E-4   9.140524E-6   -1.137476E-5   1.137476E-5   9.140524E-6   1.459227E-5   -5.121535E+1   3.878465E+1   
4.147010E+2   1.000325E+2   1.000325E+2   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   2.918106E-2   -1.967716E-2   3.085662E-5   -8.718847E-6   8.718847E-6   3.085662E-5   3.206477E-5   -1.577817E+1   7.422183E+1   
4.405120E+2   9.998681E+1   9.998681E+1   1.999000E+3   1.999000E+3   9.000000E+1   1.999000E+3   1.999000E+3   4.342853E-2   -4.094779E-2   5.351840E-5   -5.350581E-6   5.350581E-6   5.351840E-5   5.378521E-5   -5.709258E+0   8.429074E+1   
4.742980E+2   1.000022E+2   1.000022E+2   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   4.637685E-2   -4.316344E-2   5.678423E-5   -6.082721E-6   6.082721E-6   5.678423E-5   5.710909E-5   -6.114204E+0   8.388580E+1   
4.965750E+2   1.000318E+2   1.000318E+2   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   4.612280E-2   -4.448818E-2   5.748995E-5   -5.028739E-6   5.028739E-6   5.748995E-5   5.770947E-5   -4.999031E+0   8.500097E+1   
5.188670E+2   9.998211E+1   9.998211E+1   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   4.896992E-2   -4.596636E-2   6.021290E-5   -6.168166E-6   6.168166E-6   6.021290E-5   6.052800E-5   -5.848936E+0   8.415106E+1   
5.411200E+2   9.999609E+1   9.999609E+1   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   4.817103E-2   -4.775928E-2   6.088670E-5   -4.405120E-6   4.405120E-6   6.088670E-5   6.104584E-5   -4.138109E+0   8.586189E+1   
5.633730E+2   1.000690E+2   1.000690E+2   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   5.197836E-2   -4.944181E-2   6.433638E-5   -6.121151E-6   6.121151E-6   6.433638E-5   6.462692E-5   -5.434927E+0   8.456507E+1   
5.856850E+2   1.000059E+2   1.000059E+2   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   5.150162E-2   -5.165748E-2   6.548468E-5   -4.319995E-6   4.319995E-6   6.548468E-5   6.562702E-5   -3.774308E+0   8.622569E+1   
6.079350E+2   9.998708E+1   9.998708E+1   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   5.416581E-2   -5.375778E-2   6.849971E-5   -4.917396E-6   4.917396E-6   6.849971E-5   6.867598E-5   -4.106055E+0   8.589395E+1   
6.301770E+2   9.997289E+1   9.997289E+1   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   5.535617E-2   -5.509418E-2   7.010603E-5   -4.924121E-6   4.924121E-6   7.010603E-5   7.027875E-5   -4.017754E+0   8.598225E+1   
6.523990E+2   1.000019E+2   1.000019E+2   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   5.505920E-2   -5.676618E-2   7.101138E-5   -3.611365E-6   3.611365E-6   7.101138E-5   7.110316E-5   -2.911334E+0   8.708867E+1   
6.746220E+2   9.999789E+1   9.999789E+1   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   5.810749E-2   -5.781910E-2   7.358173E-5   -5.177613E-6   5.177613E-6   7.358173E-5   7.376367E-5   -4.025010E+0   8.597499E+1   
6.968940E+2   9.996520E+1   9.996520E+1   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   6.007650E-2   -6.087107E-2   7.678678E-5   -4.638656E-6   4.638656E-6   7.678678E-5   7.692676E-5   -3.457012E+0   8.654299E+1   
7.191290E+2   9.998849E+1   9.998849E+1   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   6.016115E-2   -6.272838E-2   7.804877E-5   -3.487012E-6   3.487012E-6   7.804877E-5   7.812663E-5   -2.558122E+0   8.744188E+1   
7.413650E+2   1.000398E+2   1.000398E+2   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   6.094716E-2   -6.505081E-2   8.004729E-5   -2.550031E-6   2.550031E-6   8.004729E-5   8.008790E-5   -1.824629E+0   8.817537E+1   
7.636460E+2   1.000137E+2   1.000137E+2   1.298000E+3   1.298000E+3   9.000000E+1   1.299000E+3   1.299000E+3   6.329963E-2   -6.679340E-2   8.263662E-5   -3.150735E-6   3.150735E-6   8.263662E-5   8.269666E-5   -2.183492E+0   8.781651E+1   
7.858800E+2   1.000170E+2   1.000170E+2   1.248000E+3   1.248000E+3   9.000000E+1   1.249000E+3   1.249000E+3   6.383224E-2   -6.891763E-2   8.434939E-5   -2.155908E-6   2.155908E-6   8.434939E-5   8.437694E-5   -1.464119E+0   8.853588E+1   
8.081060E+2   1.000078E+2   1.000078E+2   1.198000E+3   1.198000E+3   9.000000E+1   1.198000E+3   1.198000E+3   6.556377E-2   -7.080256E-2   8.664754E-5   -2.204288E-6   2.204288E-6   8.664754E-5   8.667558E-5   -1.457274E+0   8.854273E+1   
8.301860E+2   1.000344E+2   1.000344E+2   1.148000E+3   1.148000E+3   9.000000E+1   1.149000E+3   1.149000E+3   6.812550E-2   -7.221933E-2   8.915405E-5   -3.172773E-6   3.172773E-6   8.915405E-5   8.921049E-5   -2.038156E+0   8.796184E+1   
8.524170E+2   1.000209E+2   1.000209E+2   1.098000E+3   1.098000E+3   9.000000E+1   1.099000E+3   1.099000E+3   6.906733E-2   -7.432392E-2   9.110703E-5   -2.493468E-6   2.493468E-6   9.110703E-5   9.114115E-5   -1.567711E+0   8.843229E+1   
8.747560E+2   1.000119E+2   1.000119E+2   1.048000E+3   1.048000E+3   9.000000E+1   1.049000E+3   1.049000E+3   6.922258E-2   -7.526885E-2   9.181844E-5   -1.990526E-6   1.990526E-6   9.181844E-5   9.184001E-5   -1.241917E+0   8.875808E+1   
8.968910E+2   1.000445E+2   1.000445E+2   9.980000E+2   9.980000E+2   9.000000E+1   9.990000E+2   9.990000E+2   6.968767E-2   -7.646903E-2   9.288764E-5   -1.549878E-6   1.549878E-6   9.288764E-5   9.290057E-5   -9.559206E-1   8.904408E+1   
9.187740E+2   1.000053E+2   1.000053E+2   9.480000E+2   9.480000E+2   9.000000E+1   9.480000E+2   9.480000E+2   7.204016E-2   -8.039167E-2   9.689684E-5   -7.253402E-7   7.253402E-7   9.689684E-5   9.689956E-5   -4.288907E-1   8.957111E+1   
9.406010E+2   9.997451E+1   9.997451E+1   8.970000E+2   8.970000E+2   9.000000E+1   8.980000E+2   8.980000E+2   7.350726E-2   -7.991307E-2   9.749216E-5   -2.123345E-6   2.123345E-6   9.749216E-5   9.751528E-5   -1.247685E+0   8.875232E+1   
9.624830E+2   1.000588E+2   1.000588E+2   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   7.501605E-2   -8.266316E-2   1.002161E-4   -1.441362E-6   1.441362E-6   1.002161E-4   1.002264E-4   -8.240025E-1   8.917600E+1   
9.843320E+2   1.000783E+2   1.000783E+2   7.980000E+2   7.980000E+2   9.000000E+1   7.980000E+2   7.980000E+2   7.513754E-2   -8.495060E-2   1.017810E-4   -3.575713E-8   3.575713E-8   1.017810E-4   1.017810E-4   -2.012884E-2   8.997987E+1   
1.006179E+3   1.000015E+2   1.000015E+2   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   7.628617E-2   -8.663797E-2   1.035901E-4   2.178334E-7   -2.178334E-7   1.035901E-4   1.035903E-4   1.204837E-1   9.012048E+1   
1.028055E+3   9.999450E+1   9.999450E+1   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   7.819870E-2   -8.913709E-2   1.064001E-4   4.371235E-7   -4.371235E-7   1.064001E-4   1.064010E-4   2.353868E-1   9.023539E+1   
1.049933E+3   1.000118E+2   1.000118E+2   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   7.889208E-2   -9.026794E-2   1.075653E-4   6.635973E-7   -6.635973E-7   1.075653E-4   1.075674E-4   3.534675E-1   9.035347E+1   
1.071808E+3   1.000129E+2   1.000129E+2   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   8.060397E-2   -9.257506E-2   1.101263E-4   9.057583E-7   -9.057583E-7   1.101263E-4   1.101300E-4   4.712313E-1   9.047123E+1   
1.093681E+3   9.999291E+1   9.999291E+1   5.470000E+2   5.470000E+2   9.000000E+1   5.480000E+2   5.480000E+2   8.251406E-2   -9.397602E-2   1.122196E-4   4.089058E-7   -4.089058E-7   1.122196E-4   1.122204E-4   2.087734E-1   9.020877E+1   
1.115520E+3   1.000228E+2   1.000228E+2   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   8.279447E-2   -9.550637E-2   1.133897E-4   1.202002E-6   -1.202002E-6   1.133897E-4   1.133961E-4   6.073487E-1   9.060735E+1   
1.137355E+3   1.000580E+2   1.000580E+2   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   8.498742E-2   -9.734107E-2   1.159404E-4   7.795081E-7   -7.795081E-7   1.159404E-4   1.159430E-4   3.852139E-1   9.038521E+1   
1.159203E+3   1.000175E+2   1.000175E+2   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   8.621888E-2   -9.925548E-2   1.179486E-4   1.120262E-6   -1.120262E-6   1.179486E-4   1.179539E-4   5.441721E-1   9.054417E+1   
1.180981E+3   1.000641E+2   1.000641E+2   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   8.652200E-2   -1.014073E-1   1.195375E-4   2.302879E-6   -2.302879E-6   1.195375E-4   1.195596E-4   1.103662E+0   9.110366E+1   
1.202875E+3   1.000077E+2   1.000077E+2   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   8.909294E-2   -1.021136E-1   1.215869E-4   8.630499E-7   -8.630499E-7   1.215869E-4   1.215900E-4   4.066909E-1   9.040669E+1   
1.224656E+3   1.000341E+2   1.000341E+2   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   8.940831E-2   -1.045335E-1   1.233580E-4   2.211911E-6   -2.211911E-6   1.233580E-4   1.233778E-4   1.027251E+0   9.102725E+1   
1.246548E+3   1.000240E+2   1.000240E+2   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   9.004519E-2   -1.063179E-1   1.249138E-4   2.907385E-6   -2.907385E-6   1.249138E-4   1.249477E-4   1.333325E+0   9.133333E+1   
1.268421E+3   1.000209E+2   1.000209E+2   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   9.173876E-2   -1.077144E-1   1.268704E-4   2.567770E-6   -2.567770E-6   1.268704E-4   1.268964E-4   1.159469E+0   9.115947E+1   
1.290247E+3   1.000163E+2   1.000163E+2   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   9.226524E-2   -1.097956E-1   1.285514E-4   3.539047E-6   -3.539047E-6   1.285514E-4   1.286001E-4   1.576966E+0   9.157697E+1   
1.311985E+3   1.000680E+2   1.000680E+2   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   9.453868E-2   -1.118647E-1   1.313045E-4   3.210215E-6   -3.210215E-6   1.313045E-4   1.313437E-4   1.400524E+0   9.140052E+1   
1.345174E+3   1.000472E+2   1.000472E+2   4.600000E+1   4.600000E+1   9.000000E+1   4.700000E+1   4.700000E+1   9.569842E-2   -1.119009E-1   1.320451E-4   2.376100E-6   -2.376100E-6   1.320451E-4   1.320665E-4   1.030904E+0   9.103090E+1   
1.364196E+3   9.997170E+1   9.997170E+1   4.700000E+1   4.700000E+1   9.000000E+1   4.700000E+1   4.700000E+1   9.419877E-2   -1.114529E-1   1.308262E-4   3.192448E-6   -3.192448E-6   1.308262E-4   1.308651E-4   1.397866E+0   9.139787E+1   
1.386285E+3   1.000040E+2   1.000040E+2   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   9.425397E-2   -1.111032E-1   1.306325E-4   2.922970E-6   -2.922970E-6   1.306325E-4   1.306652E-4   1.281808E+0   9.128181E+1   
1.405343E+3   1.000276E+2   1.000276E+2   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   9.265366E-2   -1.122794E-1   1.304092E-4   4.875605E-6   -4.875605E-6   1.304092E-4   1.305003E-4   2.141118E+0   9.214112E+1   
1.427728E+3   1.000011E+2   1.000011E+2   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   9.511488E-2   -1.109958E-1   1.310949E-4   2.215995E-6   -2.215995E-6   1.310949E-4   1.311136E-4   9.684216E-1   9.096842E+1   
1.446766E+3   1.000070E+2   1.000070E+2   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   9.515476E-2   -1.117922E-1   1.316382E-4   2.707195E-6   -2.707195E-6   1.316382E-4   1.316661E-4   1.178145E+0   9.117815E+1   
1.469196E+3   1.000554E+2   1.000554E+2   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   9.388583E-2   -1.120567E-1   1.310260E-4   3.818637E-6   -3.818637E-6   1.310260E-4   1.310816E-4   1.669363E+0   9.166936E+1   
1.488222E+3   1.000143E+2   1.000143E+2   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   9.428957E-2   -1.112191E-1   1.307301E-4   2.972445E-6   -2.972445E-6   1.307301E-4   1.307639E-4   1.302525E+0   9.130253E+1   
1.510671E+3   1.000593E+2   1.000593E+2   3.100000E+1   3.100000E+1   9.000000E+1   3.100000E+1   3.100000E+1   9.523025E-2   -1.127200E-1   1.322891E-4   3.257887E-6   -3.257887E-6   1.322891E-4   1.323292E-4   1.410739E+0   9.141074E+1   
1.532093E+3   1.000691E+2   1.000691E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   9.504061E-2   -1.126930E-1   1.321543E-4   3.380505E-6   -3.380505E-6   1.321543E-4   1.321975E-4   1.465306E+0   9.146531E+1   
1.551202E+3   1.000510E+2   1.000510E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   9.487247E-2   -1.116591E-1   1.313770E-4   2.828929E-6   -2.828929E-6   1.313770E-4   1.314074E-4   1.233554E+0   9.123355E+1   
1.573610E+3   9.999960E+1   9.999960E+1   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   9.587822E-2   -1.118297E-1   1.321099E-4   2.196569E-6   -2.196569E-6   1.321099E-4   1.321281E-4   9.525596E-1   9.095256E+1   
1.592616E+3   9.994589E+1   9.994589E+1   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   9.597085E-2   -1.118824E-1   1.322015E-4   2.162557E-6   -2.162557E-6   1.322015E-4   1.322192E-4   9.371630E-1   9.093716E+1   
1.615072E+3   1.000342E+2   1.000342E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   9.489278E-2   -1.116616E-1   1.313911E-4   2.815524E-6   -2.815524E-6   1.313911E-4   1.314213E-4   1.227579E+0   9.122758E+1   
1.634100E+3   9.999941E+1   9.999941E+1   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   9.451232E-2   -1.135943E-1   1.324147E-4   4.360517E-6   -4.360517E-6   1.324147E-4   1.324865E-4   1.886112E+0   9.188611E+1   
1.656481E+3   1.000079E+2   1.000079E+2   1.700000E+1   1.700000E+1   9.000000E+1   1.700000E+1   1.700000E+1   9.500561E-2   -1.117088E-1   1.314917E-4   2.762953E-6   -2.762953E-6   1.314917E-4   1.315207E-4   1.203744E+0   9.120374E+1   
1.677870E+3   9.995959E+1   9.995959E+1   1.500000E+1   1.500000E+1   9.000000E+1   1.500000E+1   1.500000E+1   9.466571E-2   -1.121573E-1   1.315737E-4   3.307597E-6   -3.307597E-6   1.315737E-4   1.316152E-4   1.440041E+0   9.144004E+1   
1.699253E+3   1.000370E+2   1.000370E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   9.471722E-2   -1.130163E-1   1.321650E-4   3.831093E-6   -3.831093E-6   1.321650E-4   1.322205E-4   1.660380E+0   9.166038E+1   
1.718364E+3   1.000083E+2   1.000083E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   9.592545E-2   -1.129212E-1   1.328500E-4   2.875275E-6   -2.875275E-6   1.328500E-4   1.328811E-4   1.239860E+0   9.123986E+1   
1.740450E+3   1.000144E+2   1.000144E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   9.501302E-2   -1.133606E-1   1.325720E-4   3.837350E-6   -3.837350E-6   1.325720E-4   1.326275E-4   1.657986E+0   9.165799E+1   
1.759184E+3   1.000316E+2   1.000316E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   9.553092E-2   -1.136496E-1   1.330805E-4   3.643247E-6   -3.643247E-6   1.330805E-4   1.331303E-4   1.568153E+0   9.156815E+1   
1.781186E+3   9.999630E+1   9.999630E+1   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   9.614392E-2   -1.128268E-1   1.329235E-4   2.651913E-6   -2.651913E-6   1.329235E-4   1.329500E-4   1.142937E+0   9.114294E+1   
1.799953E+3   1.000667E+2   1.000667E+2   4.000000E+0   4.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   9.630034E-2   -1.123635E-1   1.327185E-4   2.233358E-6   -2.233358E-6   1.327185E-4   1.327373E-4   9.640697E-1   9.096407E+1   
1.821989E+3   1.000682E+2   1.000682E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   9.585550E-2   -1.139742E-1   1.334925E-4   3.615375E-6   -3.615375E-6   1.334925E-4   1.335415E-4   1.551361E+0   9.155136E+1   
1.840686E+3   1.000672E+2   1.000672E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   9.582668E-2   -1.140932E-1   1.335522E-4   3.714502E-6   -3.714502E-6   1.335522E-4   1.336039E-4   1.593163E+0   9.159316E+1   
1.862752E+3   9.997430E+1   9.997430E+1   -1.000000E+0   -1.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   9.667832E-2   -1.124144E-1   1.329854E-4   1.987084E-6   -1.987084E-6   1.329854E-4   1.330002E-4   8.560569E-1   9.085606E+1   
1.884481E+3   1.000622E+2   1.000622E+2   -3.000000E+0   -3.000000E+0   9.000000E+1   -3.000000E+0   -3.000000E+0   9.683113E-2   -1.130078E-1   1.334663E-4   2.261964E-6   -2.261964E-6   1.334663E-4   1.334855E-4   9.709460E-1   9.097095E+1   
1.906236E+3   1.000237E+2   1.000237E+2   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   9.502831E-2   -1.131624E-1   1.324524E-4   3.696469E-6   -3.696469E-6   1.324524E-4   1.325040E-4   1.598590E+0   9.159859E+1   
1.928254E+3   9.995989E+1   9.995989E+1   -8.000000E+0   -8.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   9.651513E-2   -1.132790E-1   1.334476E-4   2.673001E-6   -2.673001E-6   1.334476E-4   1.334743E-4   1.147501E+0   9.114750E+1   
1.950332E+3   1.000426E+2   1.000426E+2   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   9.535048E-2   -1.137171E-1   1.330128E-4   3.820837E-6   -3.820837E-6   1.330128E-4   1.330677E-4   1.645387E+0   9.164539E+1   
1.972602E+3   1.000498E+2   1.000498E+2   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   9.764479E-2   -1.138655E-1   1.345280E-4   2.220954E-6   -2.220954E-6   1.345280E-4   1.345463E-4   9.458232E-1   9.094582E+1   
1.994882E+3   1.000414E+2   1.000414E+2   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   9.611261E-2   -1.142699E-1   1.338441E-4   3.618564E-6   -3.618564E-6   1.338441E-4   1.338930E-4   1.548652E+0   9.154865E+1   
2.017124E+3   1.000410E+2   1.000410E+2   -1.500000E+1   -1.500000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   9.643658E-2   -1.136017E-1   1.336092E-4   2.942096E-6   -2.942096E-6   1.336092E-4   1.336416E-4   1.261459E+0   9.126146E+1   
2.039060E+3   1.000366E+2   1.000366E+2   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   9.507254E-2   -1.132544E-1   1.325397E-4   3.723936E-6   -3.723936E-6   1.325397E-4   1.325920E-4   1.609403E+0   9.160940E+1   
2.061256E+3   1.000289E+2   1.000289E+2   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   9.591930E-2   -1.138846E-1   1.334736E-4   3.509622E-6   -3.509622E-6   1.334736E-4   1.335197E-4   1.506217E+0   9.150622E+1   
2.083441E+3   9.996450E+1   9.996450E+1   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   9.749690E-2   -1.137680E-1   1.343730E-4   2.266563E-6   -2.266563E-6   1.343730E-4   1.343921E-4   9.663562E-1   9.096636E+1   
2.105664E+3   1.000039E+2   1.000039E+2   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   9.724899E-2   -1.146651E-1   1.348040E-4   3.036396E-6   -3.036396E-6   1.348040E-4   1.348382E-4   1.290342E+0   9.129034E+1   
2.127927E+3   1.000587E+2   1.000587E+2   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   9.721645E-2   -1.137649E-1   1.341976E-4   2.471989E-6   -2.471989E-6   1.341976E-4   1.342204E-4   1.055298E+0   9.105530E+1   
2.150185E+3   1.000007E+2   1.000007E+2   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   9.717597E-2   -1.144153E-1   1.345962E-4   2.927143E-6   -2.927143E-6   1.345962E-4   1.346280E-4   1.245849E+0   9.124585E+1   
2.172444E+3   9.998480E+1   9.998480E+1   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   9.723427E-2   -1.146865E-1   1.348089E-4   3.061329E-6   -3.061329E-6   1.348089E-4   1.348436E-4   1.300886E+0   9.130089E+1   
2.194730E+3   1.000088E+2   1.000088E+2   -3.100000E+1   -3.100000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   9.678083E-2   -1.142607E-1   1.342512E-4   3.118301E-6   -3.118301E-6   1.342512E-4   1.342874E-4   1.330591E+0   9.133059E+1   
2.216613E+3   9.995590E+1   9.995590E+1   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   9.709192E-2   -1.137576E-1   1.341159E-4   2.559272E-6   -2.559272E-6   1.341159E-4   1.341403E-4   1.093217E+0   9.109322E+1   
2.238854E+3   1.000467E+2   1.000467E+2   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   9.670416E-2   -1.135404E-1   1.337347E-4   2.704078E-6   -2.704078E-6   1.337347E-4   1.337620E-4   1.158347E+0   9.115835E+1   
2.261135E+3   1.000097E+2   1.000097E+2   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   9.700907E-2   -1.140398E-1   1.342485E-4   2.805081E-6   -2.805081E-6   1.342485E-4   1.342778E-4   1.197004E+0   9.119700E+1   
2.283387E+3   9.997820E+1   9.997820E+1   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   9.654892E-2   -1.151479E-1   1.346857E-4   3.869887E-6   -3.869887E-6   1.346857E-4   1.347413E-4   1.645811E+0   9.164581E+1   
2.305588E+3   1.000975E+2   1.000975E+2   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   9.699129E-2   -1.146540E-1   1.346375E-4   3.219764E-6   -3.219764E-6   1.346375E-4   1.346760E-4   1.369929E+0   9.136993E+1   
2.327762E+3   1.000268E+2   1.000268E+2   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   9.692686E-2   -1.152707E-1   1.349993E-4   3.670587E-6   -3.670587E-6   1.349993E-4   1.350492E-4   1.557470E+0   9.155747E+1   
2.350033E+3   9.997180E+1   9.997180E+1   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   9.723240E-2   -1.144969E-1   1.346843E-4   2.938749E-6   -2.938749E-6   1.346843E-4   1.347163E-4   1.249969E+0   9.124997E+1   
2.372292E+3   1.000655E+2   1.000655E+2   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   9.679984E-2   -1.150449E-1   1.347737E-4   3.616910E-6   -3.616910E-6   1.347737E-4   1.348222E-4   1.537273E+0   9.153727E+1   
2.394535E+3   9.998290E+1   9.998290E+1   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   9.787793E-2   -1.144258E-1   1.350370E-4   2.414777E-6   -2.414777E-6   1.350370E-4   1.350586E-4   1.024473E+0   9.102447E+1   
2.427889E+3   9.999990E+1   9.999990E+1   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   9.880017E-2   -1.167782E-1   1.371393E-4   3.270639E-6   -3.270639E-6   1.371393E-4   1.371783E-4   1.366190E+0   9.136619E+1   
2.449665E+3   1.000256E+2   1.000256E+2   -1.510000E+2   -1.510000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   9.981322E-2   -1.172139E-1   1.380494E-4   2.806167E-6   -2.806167E-6   1.380494E-4   1.380779E-4   1.164506E+0   9.116451E+1   
2.471346E+3   1.000181E+2   1.000181E+2   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   1.017393E-1   -1.201763E-1   1.411695E-4   3.318337E-6   -3.318337E-6   1.411695E-4   1.412085E-4   1.346549E+0   9.134655E+1   
2.493050E+3   1.000205E+2   1.000205E+2   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   1.006054E-1   -1.210107E-1   1.410120E-4   4.702545E-6   -4.702545E-6   1.410120E-4   1.410904E-4   1.910023E+0   9.191002E+1   
2.514789E+3   1.000140E+2   1.000140E+2   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   1.022038E-1   -1.232356E-1   1.434492E-4   4.974895E-6   -4.974895E-6   1.434492E-4   1.435354E-4   1.986252E+0   9.198625E+1   
2.536485E+3   1.000423E+2   1.000423E+2   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   1.026259E-1   -1.252997E-1   1.450545E-4   6.012102E-6   -6.012102E-6   1.450545E-4   1.451790E-4   2.373391E+0   9.237339E+1   
2.558227E+3   9.995901E+1   9.995901E+1   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   1.056650E-1   -1.269723E-1   1.480228E-4   4.857821E-6   -4.857821E-6   1.480228E-4   1.481025E-4   1.879662E+0   9.187966E+1   
2.580666E+3   1.000458E+2   1.000458E+2   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   1.064393E-1   -1.276418E-1   1.489375E-4   4.722746E-6   -4.722746E-6   1.489375E-4   1.490124E-4   1.816217E+0   9.181622E+1   
2.602352E+3   1.000114E+2   1.000114E+2   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   1.073836E-1   -1.290598E-1   1.504448E-4   4.951359E-6   -4.951359E-6   1.504448E-4   1.505263E-4   1.885007E+0   9.188501E+1   
2.624089E+3   1.000253E+2   1.000253E+2   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   1.086071E-1   -1.309238E-1   1.524153E-4   5.265079E-6   -5.265079E-6   1.524153E-4   1.525062E-4   1.978455E+0   9.197846E+1   
2.645793E+3   9.999771E+1   9.999771E+1   -6.000000E+2   -6.000000E+2   9.000000E+1   -5.990000E+2   -5.990000E+2   1.109283E-1   -1.316920E-1   1.543507E-4   4.050497E-6   -4.050497E-6   1.543507E-4   1.544038E-4   1.503220E+0   9.150322E+1   
2.667478E+3   1.000502E+2   1.000502E+2   -6.500000E+2   -6.500000E+2   9.000000E+1   -6.490000E+2   -6.490000E+2   1.115634E-1   -1.341421E-1   1.563390E-4   5.182558E-6   -5.182558E-6   1.563390E-4   1.564249E-4   1.898630E+0   9.189863E+1   
2.689150E+3   1.000348E+2   1.000348E+2   -7.010000E+2   -7.010000E+2   9.000000E+1   -7.000000E+2   -7.000000E+2   1.115842E-1   -1.353343E-1   1.571284E-4   5.946571E-6   -5.946571E-6   1.571284E-4   1.572409E-4   2.167342E+0   9.216734E+1   
2.710837E+3   1.000193E+2   1.000193E+2   -7.510000E+2   -7.510000E+2   9.000000E+1   -7.490000E+2   -7.490000E+2   1.124273E-1   -1.372616E-1   1.589048E-4   6.583000E-6   -6.583000E-6   1.589048E-4   1.590411E-4   2.372254E+0   9.237225E+1   
2.732567E+3   1.000705E+2   1.000705E+2   -8.010000E+2   -8.010000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   1.139508E-1   -1.389011E-1   1.609145E-4   6.528000E-6   -6.528000E-6   1.609145E-4   1.610469E-4   2.323108E+0   9.232311E+1   
2.754283E+3   1.000337E+2   1.000337E+2   -8.500000E+2   -8.500000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   1.147853E-1   -1.397607E-1   1.619903E-4   6.472805E-6   -6.472805E-6   1.619903E-4   1.621196E-4   2.288206E+0   9.228821E+1   
2.775908E+3   1.000298E+2   1.000298E+2   -9.000000E+2   -9.000000E+2   9.000000E+1   -9.000000E+2   -9.000000E+2   1.167206E-1   -1.420144E-1   1.646546E-4   6.514843E-6   -6.514843E-6   1.646546E-4   1.647834E-4   2.265825E+0   9.226582E+1   
2.797538E+3   1.000514E+2   1.000514E+2   -9.510000E+2   -9.510000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   1.177330E-1   -1.435631E-1   1.662891E-4   6.778509E-6   -6.778509E-6   1.662891E-4   1.664272E-4   2.334278E+0   9.233428E+1   
2.819282E+3   1.000007E+2   1.000007E+2   -1.000000E+3   -1.000000E+3   9.000000E+1   -1.000000E+3   -1.000000E+3   1.194522E-1   -1.455419E-1   1.686409E-4   6.800586E-6   -6.800586E-6   1.686409E-4   1.687779E-4   2.309250E+0   9.230925E+1   
2.841415E+3   1.000296E+2   1.000296E+2   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.049000E+3   -1.049000E+3   1.194596E-1   -1.475403E-1   1.699470E-4   8.101666E-6   -8.101666E-6   1.699470E-4   1.701400E-4   2.729323E+0   9.272932E+1   
2.863299E+3   1.000057E+2   1.000057E+2   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   1.205659E-1   -1.496063E-1   1.719765E-4   8.634054E-6   -8.634054E-6   1.719765E-4   1.721931E-4   2.874113E+0   9.287411E+1   
2.885176E+3   1.000616E+2   1.000616E+2   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.149000E+3   -1.149000E+3   1.232779E-1   -1.510746E-1   1.746095E-4   7.588089E-6   -7.588089E-6   1.746095E-4   1.747743E-4   2.488365E+0   9.248837E+1   
2.907783E+3   9.999029E+1   9.999029E+1   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   1.233007E-1   -1.526435E-1   1.756453E-4   8.597023E-6   -8.597023E-6   1.756453E-4   1.758556E-4   2.802126E+0   9.280213E+1   
2.929826E+3   1.000075E+2   1.000075E+2   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   1.241854E-1   -1.540265E-1   1.770931E-4   8.846800E-6   -8.846800E-6   1.770931E-4   1.773139E-4   2.859870E+0   9.285987E+1   
2.951675E+3   1.000317E+2   1.000317E+2   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   1.257648E-1   -1.550414E-1   1.787305E-4   8.342137E-6   -8.342137E-6   1.787305E-4   1.789251E-4   2.672306E+0   9.267231E+1   
2.974286E+3   1.000253E+2   1.000253E+2   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   1.255157E-1   -1.576215E-1   1.802569E-4   1.021319E-5   -1.021319E-5   1.802569E-4   1.805460E-4   3.242857E+0   9.324286E+1   
2.996425E+3   9.998889E+1   9.998889E+1   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   1.274767E-1   -1.586045E-1   1.821095E-4   9.405402E-6   -9.405402E-6   1.821095E-4   1.823522E-4   2.956526E+0   9.295653E+1   
3.018563E+3   1.000339E+2   1.000339E+2   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   1.282860E-1   -1.609017E-1   1.841060E-4   1.030870E-5   -1.030870E-5   1.841060E-4   1.843944E-4   3.204831E+0   9.320483E+1   
3.040951E+3   9.998980E+1   9.998980E+1   -1.500000E+3   -1.500000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   1.284811E-1   -1.627100E-1   1.854043E-4   1.134656E-5   -1.134656E-5   1.854043E-4   1.857512E-4   3.502078E+0   9.350208E+1   
3.063080E+3   1.000459E+2   1.000459E+2   -1.549000E+3   -1.549000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   1.300869E-1   -1.621915E-1   1.860594E-4   9.819928E-6   -9.819928E-6   1.860594E-4   1.863184E-4   3.021180E+0   9.302118E+1   
3.085206E+3   1.000323E+2   1.000323E+2   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.598000E+3   -1.598000E+3   1.313337E-1   -1.637279E-1   1.878309E-4   9.902214E-6   -9.902214E-6   1.878309E-4   1.880917E-4   3.017769E+0   9.301777E+1   
3.108077E+3   1.000535E+2   1.000535E+2   -1.649000E+3   -1.649000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   1.342697E-1   -1.667455E-1   1.916114E-4   9.703470E-6   -9.703470E-6   1.916114E-4   1.918570E-4   2.899062E+0   9.289906E+1   
3.130196E+3   1.000308E+2   1.000308E+2   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.698000E+3   -1.698000E+3   1.333401E-1   -1.690183E-1   1.925169E-4   1.187687E-5   -1.187687E-5   1.925169E-4   1.928829E-4   3.530253E+0   9.353025E+1   
3.152325E+3   1.000388E+2   1.000388E+2   -1.749000E+3   -1.749000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   1.332512E-1   -1.694324E-1   1.927316E-4   1.221344E-5   -1.221344E-5   1.927316E-4   1.931182E-4   3.625996E+0   9.362600E+1   
3.175558E+3   9.999249E+1   9.999249E+1   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.799000E+3   -1.799000E+3   1.342071E-1   -1.712726E-1   1.945211E-4   1.270942E-5   -1.270942E-5   1.945211E-4   1.949359E-4   3.738220E+0   9.373822E+1   
3.197681E+3   9.995779E+1   9.995779E+1   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.848000E+3   -1.848000E+3   1.348152E-1   -1.721592E-1   1.954745E-4   1.283934E-5   -1.283934E-5   1.954745E-4   1.958957E-4   3.757956E+0   9.375796E+1   
3.220306E+3   1.000412E+2   1.000412E+2   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.898000E+3   -1.898000E+3   1.375027E-1   -1.728605E-1   1.975928E-4   1.131007E-5   -1.131007E-5   1.975928E-4   1.979162E-4   3.275995E+0   9.327600E+1   
3.243190E+3   1.000374E+2   1.000374E+2   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.948000E+3   -1.948000E+3   1.373395E-1   -1.760211E-1   1.995504E-4   1.349708E-5   -1.349708E-5   1.995504E-4   2.000063E-4   3.869448E+0   9.386945E+1   
3.265488E+3   9.999670E+1   9.999670E+1   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   1.385667E-1   -1.783926E-1   2.018536E-4   1.413985E-5   -1.413985E-5   2.018536E-4   2.023482E-4   4.007026E+0   9.400703E+1   
3.302538E+3   1.000564E+2   1.000564E+2   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   1.522772E-1   -1.965751E-1   2.221722E-4   1.588629E-5   -1.588629E-5   2.221722E-4   2.227394E-4   4.089942E+0   9.408994E+1   
3.329052E+3   9.999691E+1   9.999691E+1   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.625400E-1   -2.133585E-1   2.394480E-4   1.926810E-5   -1.926810E-5   2.394480E-4   2.402220E-4   4.600613E+0   9.460061E+1   
3.354184E+3   1.000481E+2   1.000481E+2   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.755419E-1   -2.330650E-1   2.603210E-4   2.253507E-5   -2.253507E-5   2.603210E-4   2.612945E-4   4.947559E+0   9.494756E+1   
3.379791E+3   1.000495E+2   1.000495E+2   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   1.865462E-1   -2.478525E-1   2.767552E-4   2.406361E-5   -2.406361E-5   2.767552E-4   2.777994E-4   4.969316E+0   9.496932E+1   
3.405592E+3   1.000197E+2   1.000197E+2   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   1.922075E-1   -2.603107E-1   2.883692E-4   2.802119E-5   -2.802119E-5   2.883692E-4   2.897275E-4   5.550076E+0   9.555008E+1   
3.430318E+3   9.999951E+1   9.999951E+1   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   1.936108E-1   -2.665024E-1   2.932694E-4   3.103115E-5   -3.103115E-5   2.932694E-4   2.949066E-4   6.040053E+0   9.604005E+1   
3.455491E+3   9.996539E+1   9.996539E+1   -5.500000E+3   -5.500000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   1.852839E-1   -2.572863E-1   2.821191E-4   3.116479E-5   -3.116479E-5   2.821191E-4   2.838352E-4   6.303722E+0   9.630372E+1   
3.481641E+3   1.000076E+2   1.000076E+2   -6.000000E+3   -6.000000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   1.751007E-1   -2.441053E-1   2.672386E-4   3.007919E-5   -3.007919E-5   2.672386E-4   2.689261E-4   6.421930E+0   9.642193E+1   
3.506379E+3   9.998889E+1   9.998889E+1   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   1.594482E-1   -2.282686E-1   2.472472E-4   3.130275E-5   -3.130275E-5   2.472472E-4   2.492209E-4   7.215546E+0   9.721555E+1   
3.531040E+3   1.000255E+2   1.000255E+2   -7.000000E+3   -7.000000E+3   9.000000E+1   -7.000000E+3   -7.000000E+3   1.537062E-1   -2.222064E-1   2.397490E-4   3.158636E-5   -3.158636E-5   2.397490E-4   2.418208E-4   7.505356E+0   9.750536E+1   
3.556240E+3   1.000099E+2   1.000099E+2   -7.500000E+3   -7.500000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.521766E-1   -2.203816E-1   2.376149E-4   3.152473E-5   -3.152473E-5   2.376149E-4   2.396970E-4   7.557385E+0   9.755738E+1   
3.581433E+3   1.000028E+2   1.000028E+2   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.569656E-1   -2.296240E-1   2.465952E-4   3.402504E-5   -3.402504E-5   2.465952E-4   2.489315E-4   7.856031E+0   9.785603E+1   
3.607123E+3   9.995849E+1   9.995849E+1   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.649005E-1   -2.399776E-1   2.582441E-4   3.492507E-5   -3.492507E-5   2.582441E-4   2.605950E-4   7.701983E+0   9.770198E+1   
3.632818E+3   1.000102E+2   1.000102E+2   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.785607E-1   -2.577196E-1   2.782446E-4   3.642070E-5   -3.642070E-5   2.782446E-4   2.806181E-4   7.457308E+0   9.745731E+1   
3.658522E+3   1.000509E+2   1.000509E+2   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.919325E-1   -2.759994E-1   2.984172E-4   3.848138E-5   -3.848138E-5   2.984172E-4   3.008881E-4   7.347836E+0   9.734784E+1   
3.683695E+3   1.000827E+2   1.000827E+2   -9.999000E+3   -9.999000E+3   9.000000E+1   -9.998000E+3   -9.998000E+3   2.062090E-1   -2.966072E-1   3.206652E-4   4.139485E-5   -4.139485E-5   3.206652E-4   3.233260E-4   7.355666E+0   9.735567E+1   
3.720176E+3   9.997439E+1   9.997439E+1   -9.500000E+3   -9.500000E+3   9.000000E+1   -9.499000E+3   -9.499000E+3   1.815980E-1   -2.665728E-1   2.858885E-4   3.996227E-5   -3.996227E-5   2.858885E-4   2.886680E-4   7.957400E+0   9.795740E+1   
3.744865E+3   1.000344E+2   1.000344E+2   -9.000000E+3   -9.000000E+3   9.000000E+1   -8.999000E+3   -8.999000E+3   1.639635E-1   -2.439286E-1   2.602380E-4   3.820107E-5   -3.820107E-5   2.602380E-4   2.630269E-4   8.350968E+0   9.835097E+1   
3.769539E+3   1.000376E+2   1.000376E+2   -8.500000E+3   -8.500000E+3   9.000000E+1   -8.499000E+3   -8.499000E+3   1.464107E-1   -2.208037E-1   2.343251E-4   3.606532E-5   -3.606532E-5   2.343251E-4   2.370843E-4   8.749818E+0   9.874982E+1   
3.794229E+3   1.000410E+2   1.000410E+2   -7.999000E+3   -7.999000E+3   9.000000E+1   -7.998000E+3   -7.998000E+3   1.323977E-1   -1.998504E-1   2.120149E-4   3.273112E-5   -3.273112E-5   2.120149E-4   2.145265E-4   8.776109E+0   9.877611E+1   
3.818952E+3   1.001198E+2   1.001198E+2   -7.499000E+3   -7.499000E+3   9.000000E+1   -7.499000E+3   -7.499000E+3   1.165310E-1   -1.801671E-1   1.893858E-4   3.159824E-5   -3.159824E-5   1.893858E-4   1.920037E-4   9.472312E+0   9.947231E+1   
3.843657E+3   1.000757E+2   1.000757E+2   -7.000000E+3   -7.000000E+3   9.000000E+1   -6.999000E+3   -6.999000E+3   9.940575E-2   -1.578437E-1   1.642592E-4   2.967015E-5   -2.967015E-5   1.642592E-4   1.669173E-4   1.023894E+1   1.002389E+2   
3.868351E+3   9.998641E+1   9.998641E+1   -6.500000E+3   -6.500000E+3   9.000000E+1   -6.499000E+3   -6.499000E+3   8.664717E-2   -1.405682E-1   1.451199E-4   2.781256E-5   -2.781256E-5   1.451199E-4   1.477610E-4   1.084931E+1   1.008493E+2   
3.892498E+3   1.000509E+2   1.000509E+2   -5.999000E+3   -5.999000E+3   9.000000E+1   -5.999000E+3   -5.999000E+3   6.778188E-2   -1.185392E-1   1.191093E-4   2.736401E-5   -2.736401E-5   1.191093E-4   1.222121E-4   1.293855E+1   1.029385E+2   
3.917291E+3   1.000520E+2   1.000520E+2   -5.499000E+3   -5.499000E+3   9.000000E+1   -5.499000E+3   -5.499000E+3   5.847010E-2   -1.018270E-1   1.024678E-4   2.332532E-5   -2.332532E-5   1.024678E-4   1.050891E-4   1.282403E+1   1.028240E+2   
3.942499E+3   1.000392E+2   1.000392E+2   -5.000000E+3   -5.000000E+3   9.000000E+1   -4.999000E+3   -4.999000E+3   4.617069E-2   -8.275580E-2   8.244285E-5   1.995413E-5   -1.995413E-5   8.244285E-5   8.482330E-5   1.360598E+1   1.036060E+2   
3.966757E+3   1.000243E+2   1.000243E+2   -4.500000E+3   -4.500000E+3   9.000000E+1   -4.499000E+3   -4.499000E+3   3.510215E-2   -6.649704E-2   6.501061E-5   1.751124E-5   -1.751124E-5   6.501061E-5   6.732773E-5   1.507538E+1   1.050754E+2   
3.991426E+3   1.000457E+2   1.000457E+2   -3.999000E+3   -3.999000E+3   9.000000E+1   -3.998000E+3   -3.998000E+3   2.437727E-2   -4.832442E-2   4.654435E-5   1.356296E-5   -1.356296E-5   4.654435E-5   4.848021E-5   1.624605E+1   1.062460E+2   
4.016207E+3   9.997051E+1   9.997051E+1   -3.500000E+3   -3.500000E+3   9.000000E+1   -3.499000E+3   -3.499000E+3   1.194902E-2   -3.072605E-2   2.739899E-5   1.124996E-5   -1.124996E-5   2.739899E-5   2.961868E-5   2.232293E+1   1.123229E+2   
4.040385E+3   9.997799E+1   9.997799E+1   -3.000000E+3   -3.000000E+3   9.000000E+1   -2.999000E+3   -2.999000E+3   1.816213E-4   -1.414935E-2   9.327610E-6   9.116115E-6   -9.116115E-6   9.327610E-6   1.304254E-5   4.434301E+1   1.343430E+2   
4.065142E+3   9.999310E+1   9.999310E+1   -2.500000E+3   -2.500000E+3   9.000000E+1   -2.499000E+3   -2.499000E+3   -1.452426E-2   4.631980E-3   -1.199634E-5   7.714336E-6   -7.714336E-6   -1.199634E-5   1.426265E-5   1.472566E+2   2.372566E+2   
4.089788E+3   1.000304E+2   1.000304E+2   -1.999000E+3   -1.999000E+3   9.000000E+1   -1.998000E+3   -1.998000E+3   -2.554001E-2   2.264204E-2   -3.053655E-5   4.087459E-6   -4.087459E-6   -3.053655E-5   3.080890E-5   1.723760E+2   2.623760E+2   
4.123478E+3   1.000287E+2   1.000287E+2   -1.949000E+3   -1.949000E+3   9.000000E+1   -1.949000E+3   -1.949000E+3   -2.262484E-2   2.374895E-2   -2.945518E-5   1.207645E-6   -1.207645E-6   -2.945518E-5   2.947992E-5   1.776522E+2   2.676522E+2   
4.145510E+3   1.000098E+2   1.000098E+2   -1.899000E+3   -1.899000E+3   9.000000E+1   -1.899000E+3   -1.899000E+3   -2.281015E-2   2.568669E-2   -3.083177E-5   7.786289E-8   -7.786289E-8   -3.083177E-5   3.083187E-5   1.798553E+2   2.698553E+2   
4.167600E+3   1.000319E+2   1.000319E+2   -1.849000E+3   -1.849000E+3   9.000000E+1   -1.849000E+3   -1.849000E+3   -2.387842E-2   2.772440E-2   -3.281936E-5   -4.642128E-7   4.642128E-7   -3.281936E-5   3.282265E-5   -1.791896E+2   -8.918964E+1   
4.189382E+3   1.000154E+2   1.000154E+2   -1.799000E+3   -1.799000E+3   9.000000E+1   -1.798000E+3   -1.798000E+3   -2.576583E-2   2.975474E-2   -3.530859E-5   -3.956029E-7   3.956029E-7   -3.530859E-5   3.531081E-5   -1.793581E+2   -8.935808E+1   
4.211466E+3   9.997479E+1   9.997479E+1   -1.750000E+3   -1.750000E+3   9.000000E+1   -1.749000E+3   -1.749000E+3   -2.673713E-2   3.014684E-2   -3.616446E-5   6.645901E-8   -6.645901E-8   -3.616446E-5   3.616452E-5   1.798947E+2   2.698947E+2   
4.233497E+3   1.000300E+2   1.000300E+2   -1.699000E+3   -1.699000E+3   9.000000E+1   -1.699000E+3   -1.699000E+3   -2.802997E-2   3.165504E-2   -3.794603E-5   3.666539E-8   -3.666539E-8   -3.794603E-5   3.794605E-5   1.799446E+2   2.699446E+2   
4.255623E+3   1.000387E+2   1.000387E+2   -1.650000E+3   -1.650000E+3   9.000000E+1   -1.649000E+3   -1.649000E+3   -2.981858E-2   3.484445E-2   -4.112906E-5   -7.255733E-7   7.255733E-7   -4.112906E-5   4.113546E-5   -1.789893E+2   -8.898933E+1   
4.277385E+3   1.000778E+2   1.000778E+2   -1.599000E+3   -1.599000E+3   9.000000E+1   -1.599000E+3   -1.599000E+3   -3.055427E-2   3.605874E-2   -4.237476E-5   -9.752965E-7   9.752965E-7   -4.237476E-5   4.238598E-5   -1.786815E+2   -8.868151E+1   
4.299451E+3   1.000336E+2   1.000336E+2   -1.550000E+3   -1.550000E+3   9.000000E+1   -1.549000E+3   -1.549000E+3   -3.228887E-2   3.758042E-2   -4.443822E-5   -6.871686E-7   6.871686E-7   -4.443822E-5   4.444353E-5   -1.791141E+2   -8.911408E+1   
4.321320E+3   1.000439E+2   1.000439E+2   -1.499000E+3   -1.499000E+3   9.000000E+1   -1.499000E+3   -1.499000E+3   -3.361483E-2   3.997465E-2   -4.681733E-5   -1.271725E-6   1.271725E-6   -4.681733E-5   4.683460E-5   -1.784440E+2   -8.844403E+1   
4.343433E+3   9.998290E+1   9.998290E+1   -1.450000E+3   -1.450000E+3   9.000000E+1   -1.449000E+3   -1.449000E+3   -3.524940E-2   4.159327E-2   -4.888208E-5   -1.120949E-6   1.120949E-6   -4.888208E-5   4.889493E-5   -1.786863E+2   -8.868634E+1   
4.365542E+3   1.000293E+2   1.000293E+2   -1.400000E+3   -1.400000E+3   9.000000E+1   -1.399000E+3   -1.399000E+3   -3.605750E-2   4.286587E-2   -5.021052E-5   -1.355250E-6   1.355250E-6   -5.021052E-5   5.022881E-5   -1.784539E+2   -8.845388E+1   
4.387434E+3   1.000586E+2   1.000586E+2   -1.350000E+3   -1.350000E+3   9.000000E+1   -1.349000E+3   -1.349000E+3   -3.740676E-2   4.506067E-2   -5.247415E-5   -1.792188E-6   1.792188E-6   -5.247415E-5   5.250474E-5   -1.780439E+2   -8.804390E+1   
4.409551E+3   9.998580E+1   9.998580E+1   -1.300000E+3   -1.300000E+3   9.000000E+1   -1.299000E+3   -1.299000E+3   -3.955433E-2   4.808881E-2   -5.577407E-5   -2.183495E-6   2.183495E-6   -5.577407E-5   5.581679E-5   -1.777581E+2   -8.775808E+1   
4.431599E+3   1.000357E+2   1.000357E+2   -1.250000E+3   -1.250000E+3   9.000000E+1   -1.249000E+3   -1.249000E+3   -3.982368E-2   4.796056E-2   -5.585706E-5   -1.900427E-6   1.900427E-6   -5.585706E-5   5.588938E-5   -1.780514E+2   -8.805137E+1   
4.453470E+3   1.000527E+2   1.000527E+2   -1.200000E+3   -1.200000E+3   9.000000E+1   -1.199000E+3   -1.199000E+3   -4.058084E-2   5.136844E-2   -5.854470E-5   -3.568387E-6   3.568387E-6   -5.854470E-5   5.865334E-5   -1.765121E+2   -8.651205E+1   
4.475556E+3   1.000149E+2   1.000149E+2   -1.150000E+3   -1.150000E+3   9.000000E+1   -1.150000E+3   -1.150000E+3   -4.229584E-2   5.302147E-2   -6.068159E-5   -3.380615E-6   3.380615E-6   -6.068159E-5   6.077568E-5   -1.768113E+2   -8.681131E+1   
4.497603E+3   1.000594E+2   1.000594E+2   -1.100000E+3   -1.100000E+3   9.000000E+1   -1.099000E+3   -1.099000E+3   -4.315976E-2   5.354058E-2   -6.155380E-5   -3.081015E-6   3.081015E-6   -6.155380E-5   6.163086E-5   -1.771345E+2   -8.713451E+1   
4.519690E+3   1.000217E+2   1.000217E+2   -1.050000E+3   -1.050000E+3   9.000000E+1   -1.050000E+3   -1.050000E+3   -4.402799E-2   5.456770E-2   -6.275952E-5   -3.110353E-6   3.110353E-6   -6.275952E-5   6.283655E-5   -1.771628E+2   -8.716275E+1   
4.541678E+3   1.000530E+2   1.000530E+2   -1.000000E+3   -1.000000E+3   9.000000E+1   -9.990000E+2   -9.990000E+2   -4.463241E-2   5.704291E-2   -6.474529E-5   -4.281525E-6   4.281525E-6   -6.474529E-5   6.488670E-5   -1.762166E+2   -8.621661E+1   
4.563572E+3   1.000444E+2   1.000444E+2   -9.510000E+2   -9.510000E+2   9.000000E+1   -9.500000E+2   -9.500000E+2   -4.651308E-2   5.910823E-2   -6.725313E-5   -4.240773E-6   4.240773E-6   -6.725313E-5   6.738670E-5   -1.763919E+2   -8.639188E+1   
4.585304E+3   1.000523E+2   1.000523E+2   -9.000000E+2   -9.000000E+2   9.000000E+1   -9.000000E+2   -9.000000E+2   -4.671985E-2   6.046120E-2   -6.826214E-5   -4.972371E-6   4.972371E-6   -6.826214E-5   6.844300E-5   -1.758338E+2   -8.583380E+1   
4.607284E+3   9.999340E+1   9.999340E+1   -8.510000E+2   -8.510000E+2   9.000000E+1   -8.500000E+2   -8.500000E+2   -4.796732E-2   6.257805E-2   -7.041206E-5   -5.433641E-6   5.433641E-6   -7.041206E-5   7.062141E-5   -1.755873E+2   -8.558728E+1   
4.628922E+3   9.998019E+1   9.998019E+1   -8.000000E+2   -8.000000E+2   9.000000E+1   -7.990000E+2   -7.990000E+2   -4.854960E-2   6.348923E-2   -7.136550E-5   -5.598674E-6   5.598674E-6   -7.136550E-5   7.158477E-5   -1.755143E+2   -8.551429E+1   
4.650594E+3   9.997961E+1   9.997961E+1   -7.500000E+2   -7.500000E+2   9.000000E+1   -7.500000E+2   -7.500000E+2   -5.105492E-2   6.598285E-2   -7.453847E-5   -5.375919E-6   5.375919E-6   -7.453847E-5   7.473208E-5   -1.758748E+2   -8.587481E+1   
4.672585E+3   9.999429E+1   9.999429E+1   -7.000000E+2   -7.000000E+2   9.000000E+1   -6.990000E+2   -6.990000E+2   -5.110709E-2   6.698115E-2   -7.522091E-5   -5.989997E-6   5.989997E-6   -7.522091E-5   7.545903E-5   -1.754470E+2   -8.544703E+1   
4.694555E+3   1.000120E+2   1.000120E+2   -6.510000E+2   -6.510000E+2   9.000000E+1   -6.500000E+2   -6.500000E+2   -5.135435E-2   6.817765E-2   -7.615305E-5   -6.589352E-6   6.589352E-6   -7.615305E-5   7.643759E-5   -1.750546E+2   -8.505464E+1   
4.716144E+3   9.999529E+1   9.999529E+1   -6.000000E+2   -6.000000E+2   9.000000E+1   -6.000000E+2   -6.000000E+2   -5.452660E-2   6.972080E-2   -7.911932E-5   -5.251925E-6   5.251925E-6   -7.911932E-5   7.929343E-5   -1.762023E+2   -8.620229E+1   
4.737816E+3   9.997360E+1   9.997360E+1   -5.500000E+2   -5.500000E+2   9.000000E+1   -5.490000E+2   -5.490000E+2   -5.361666E-2   7.200826E-2   -8.004654E-5   -7.420421E-6   7.420421E-6   -8.004654E-5   8.038975E-5   -1.747037E+2   -8.470374E+1   
4.759547E+3   1.000248E+2   1.000248E+2   -5.000000E+2   -5.000000E+2   9.000000E+1   -4.990000E+2   -4.990000E+2   -5.622563E-2   7.337042E-2   -8.254669E-5   -6.381289E-6   6.381289E-6   -8.254669E-5   8.279297E-5   -1.755795E+2   -8.557953E+1   
4.781181E+3   1.000221E+2   1.000221E+2   -4.500000E+2   -4.500000E+2   9.000000E+1   -4.490000E+2   -4.490000E+2   -5.610597E-2   7.554742E-2   -8.389056E-5   -7.893054E-6   7.893054E-6   -8.389056E-5   8.426107E-5   -1.746250E+2   -8.462501E+1   
4.802876E+3   9.998290E+1   9.998290E+1   -4.000000E+2   -4.000000E+2   9.000000E+1   -3.990000E+2   -3.990000E+2   -5.736198E-2   7.671569E-2   -8.542797E-5   -7.727850E-6   7.727850E-6   -8.542797E-5   8.577679E-5   -1.748311E+2   -8.483107E+1   
4.824506E+3   1.000284E+2   1.000284E+2   -3.500000E+2   -3.500000E+2   9.000000E+1   -3.490000E+2   -3.490000E+2   -5.887569E-2   7.791707E-2   -8.714626E-5   -7.393689E-6   7.393689E-6   -8.714626E-5   8.745935E-5   -1.751505E+2   -8.515051E+1   
4.846216E+3   1.000401E+2   1.000401E+2   -3.000000E+2   -3.000000E+2   9.000000E+1   -2.990000E+2   -2.990000E+2   -5.987890E-2   7.930991E-2   -8.867364E-5   -7.562288E-6   7.562288E-6   -8.867364E-5   8.899552E-5   -1.751255E+2   -8.512548E+1   
4.867856E+3   1.000020E+2   1.000020E+2   -2.500000E+2   -2.500000E+2   9.000000E+1   -2.490000E+2   -2.490000E+2   -6.141778E-2   8.144090E-2   -9.101294E-5   -7.817267E-6   7.817267E-6   -9.101294E-5   9.134804E-5   -1.750908E+2   -8.509081E+1   
4.889542E+3   1.000583E+2   1.000583E+2   -2.000000E+2   -2.000000E+2   9.000000E+1   -1.990000E+2   -1.990000E+2   -6.232895E-2   8.263493E-2   -9.235392E-5   -7.923958E-6   7.923958E-6   -9.235392E-5   9.269324E-5   -1.750960E+2   -8.509604E+1   
4.911186E+3   1.000006E+2   1.000006E+2   -1.500000E+2   -1.500000E+2   9.000000E+1   -1.490000E+2   -1.490000E+2   -6.372486E-2   8.519603E-2   -9.488496E-5   -8.565877E-6   8.565877E-6   -9.488496E-5   9.527082E-5   -1.748415E+2   -8.484152E+1   
4.932875E+3   9.998809E+1   9.998809E+1   -1.000000E+2   -1.000000E+2   9.000000E+1   -9.900000E+1   -9.900000E+1   -6.545148E-2   8.593111E-2   -9.643118E-5   -7.769386E-6   7.769386E-6   -9.643118E-5   9.674367E-5   -1.753937E+2   -8.539367E+1   
4.954407E+3   1.000332E+2   1.000332E+2   -5.000000E+1   -5.000000E+1   9.000000E+1   -4.900000E+1   -4.900000E+1   -6.588836E-2   8.746691E-2   -9.770153E-5   -8.450318E-6   8.450318E-6   -9.770153E-5   9.806629E-5   -1.750567E+2   -8.505672E+1   
4.987431E+3   9.995559E+1   9.995559E+1   -4.800000E+1   -4.800000E+1   9.000000E+1   -4.700000E+1   -4.700000E+1   -6.577792E-2   8.727365E-2   -9.750739E-5   -8.405658E-6   8.405658E-6   -9.750739E-5   9.786903E-5   -1.750730E+2   -8.507298E+1   
5.009685E+3   1.000163E+2   1.000163E+2   -4.600000E+1   -4.600000E+1   9.000000E+1   -4.500000E+1   -4.500000E+1   -6.531588E-2   8.776512E-2   -9.754182E-5   -9.068705E-6   9.068705E-6   -9.754182E-5   9.796248E-5   -1.746883E+2   -8.468834E+1   
5.031917E+3   1.000020E+2   1.000020E+2   -4.400000E+1   -4.400000E+1   9.000000E+1   -4.300000E+1   -4.300000E+1   -6.588406E-2   8.710307E-2   -9.746192E-5   -8.215629E-6   8.215629E-6   -9.746192E-5   9.780758E-5   -1.751816E+2   -8.518160E+1   
5.054136E+3   1.000457E+2   1.000457E+2   -4.200000E+1   -4.200000E+1   9.000000E+1   -4.100000E+1   -4.100000E+1   -6.593806E-2   8.812653E-2   -9.816187E-5   -8.844797E-6   8.844797E-6   -9.816187E-5   9.855954E-5   -1.748513E+2   -8.485131E+1   
5.076409E+3   1.000085E+2   1.000085E+2   -4.000000E+1   -4.000000E+1   9.000000E+1   -3.900000E+1   -3.900000E+1   -6.544782E-2   8.653611E-2   -9.682295E-5   -8.167624E-6   8.167624E-6   -9.682295E-5   9.716684E-5   -1.751782E+2   -8.517816E+1   
5.098681E+3   1.000801E+2   1.000801E+2   -3.800000E+1   -3.800000E+1   9.000000E+1   -3.700000E+1   -3.700000E+1   -6.562882E-2   8.731476E-2   -9.744199E-5   -8.542814E-6   8.542814E-6   -9.744199E-5   9.781575E-5   -1.749896E+2   -8.498965E+1   
5.120867E+3   9.998229E+1   9.998229E+1   -3.600000E+1   -3.600000E+1   9.000000E+1   -3.500000E+1   -3.500000E+1   -6.502319E-2   8.844928E-2   -9.780645E-5   -9.732467E-6   9.732467E-6   -9.780645E-5   9.828949E-5   -1.743174E+2   -8.431735E+1   
5.143125E+3   1.000371E+2   1.000371E+2   -3.400000E+1   -3.400000E+1   9.000000E+1   -3.300000E+1   -3.300000E+1   -6.572943E-2   8.794674E-2   -9.791578E-5   -8.881565E-6   8.881565E-6   -9.791578E-5   9.831777E-5   -1.748171E+2   -8.481710E+1   
5.165395E+3   9.996780E+1   9.996780E+1   -3.200000E+1   -3.200000E+1   9.000000E+1   -3.100000E+1   -3.100000E+1   -6.675475E-2   8.884871E-2   -9.913713E-5   -8.712893E-6   8.712893E-6   -9.913713E-5   9.951927E-5   -1.749773E+2   -8.497734E+1   
5.187609E+3   9.995910E+1   9.995910E+1   -3.000000E+1   -3.000000E+1   9.000000E+1   -2.900000E+1   -2.900000E+1   -6.645838E-2   8.968013E-2   -9.949539E-5   -9.475656E-6   9.475656E-6   -9.949539E-5   9.994559E-5   -1.745597E+2   -8.455972E+1   
5.209868E+3   9.998779E+1   9.998779E+1   -2.800000E+1   -2.800000E+1   9.000000E+1   -2.700000E+1   -2.700000E+1   -6.632092E-2   8.780807E-2   -9.819117E-5   -8.353423E-6   8.353423E-6   -9.819117E-5   9.854585E-5   -1.751374E+2   -8.513738E+1   
5.232136E+3   1.000041E+2   1.000041E+2   -2.600000E+1   -2.600000E+1   9.000000E+1   -2.500000E+1   -2.500000E+1   -6.531526E-2   8.928006E-2   -9.852811E-5   -1.005959E-5   1.005959E-5   -9.852811E-5   9.904031E-5   -1.741704E+2   -8.417038E+1   
5.254343E+3   9.999209E+1   9.999209E+1   -2.400000E+1   -2.400000E+1   9.000000E+1   -2.300000E+1   -2.300000E+1   -6.575276E-2   8.870145E-2   -9.842175E-5   -9.357719E-6   9.357719E-6   -9.842175E-5   9.886560E-5   -1.745688E+2   -8.456877E+1   
5.276608E+3   1.000273E+2   1.000273E+2   -2.200000E+1   -2.200000E+1   9.000000E+1   -2.100000E+1   -2.100000E+1   -6.621847E-2   8.871494E-2   -9.871846E-5   -9.022085E-6   9.022085E-6   -9.871846E-5   9.912988E-5   -1.747781E+2   -8.477813E+1   
5.298848E+3   9.998879E+1   9.998879E+1   -2.000000E+1   -2.000000E+1   9.000000E+1   -1.900000E+1   -1.900000E+1   -6.779905E-2   8.952735E-2   -1.002248E-4   -8.384164E-6   8.384164E-6   -1.002248E-4   1.005748E-4   -1.752181E+2   -8.521813E+1   
5.321035E+3   1.000088E+2   1.000088E+2   -1.800000E+1   -1.800000E+1   9.000000E+1   -1.700000E+1   -1.700000E+1   -6.757755E-2   8.848731E-2   -9.941045E-5   -7.868051E-6   7.868051E-6   -9.941045E-5   9.972133E-5   -1.754746E+2   -8.547464E+1   
5.343297E+3   1.000108E+2   1.000108E+2   -1.600000E+1   -1.600000E+1   9.000000E+1   -1.500000E+1   -1.500000E+1   -6.616447E-2   8.874931E-2   -9.870745E-5   -9.084490E-6   9.084490E-6   -9.870745E-5   9.912461E-5   -1.747416E+2   -8.474163E+1   
5.365610E+3   1.000175E+2   1.000175E+2   -1.400000E+1   -1.400000E+1   9.000000E+1   -1.300000E+1   -1.300000E+1   -6.516432E-2   8.870331E-2   -9.805915E-5   -9.794159E-6   9.794159E-6   -9.805915E-5   9.854706E-5   -1.742962E+2   -8.429621E+1   
5.387839E+3   1.000384E+2   1.000384E+2   -1.200000E+1   -1.200000E+1   9.000000E+1   -1.100000E+1   -1.100000E+1   -6.642525E-2   8.967154E-2   -9.946932E-5   -9.494545E-6   9.494545E-6   -9.946932E-5   9.992143E-5   -1.745475E+2   -8.454752E+1   
5.409980E+3   1.000374E+2   1.000374E+2   -1.000000E+1   -1.000000E+1   9.000000E+1   -9.000000E+0   -9.000000E+0   -6.712287E-2   8.891681E-2   -9.940907E-5   -8.485141E-6   8.485141E-6   -9.940907E-5   9.977054E-5   -1.751213E+2   -8.512130E+1   
5.432120E+3   1.000496E+2   1.000496E+2   -8.000000E+0   -8.000000E+0   9.000000E+1   -7.000000E+0   -7.000000E+0   -6.615340E-2   8.927148E-2   -9.904070E-5   -9.434062E-6   9.434062E-6   -9.904070E-5   9.948900E-5   -1.745587E+2   -8.455874E+1   
5.454189E+3   1.000234E+2   1.000234E+2   -6.000000E+0   -6.000000E+0   9.000000E+1   -5.000000E+0   -5.000000E+0   -6.533430E-2   9.055818E-2   -9.937230E-5   -1.088110E-5   1.088110E-5   -9.937230E-5   9.996626E-5   -1.737511E+2   -8.375110E+1   
5.476272E+3   1.000062E+2   1.000062E+2   -4.000000E+0   -4.000000E+0   9.000000E+1   -2.000000E+0   -2.000000E+0   -6.651851E-2   8.943898E-2   -9.937551E-5   -9.273529E-6   9.273529E-6   -9.937551E-5   9.980727E-5   -1.746687E+2   -8.466871E+1   
5.498398E+3   1.000025E+2   1.000025E+2   -2.000000E+0   -2.000000E+0   9.000000E+1   -1.000000E+0   -1.000000E+0   -6.560426E-2   8.911807E-2   -9.860128E-5   -9.739930E-6   9.739930E-6   -9.860128E-5   9.908117E-5   -1.743586E+2   -8.435857E+1   
5.520443E+3   1.000587E+2   1.000587E+2   0.000000E+0   0.000000E+0   9.000000E+1   0.000000E+0   0.000000E+0   -6.594298E-2   9.005012E-2   -9.941772E-5   -1.009875E-5   1.009875E-5   -9.941772E-5   9.992931E-5   -1.741998E+2   -8.419985E+1   
5.542474E+3   1.000244E+2   1.000244E+2   0.000000E+0   0.000000E+0   9.000000E+1   1.000000E+0   1.000000E+0   -6.695354E-2   8.968627E-2   -9.980553E-5   -9.113438E-6   9.113438E-6   -9.980553E-5   1.002207E-4   -1.747827E+2   -8.478268E+1   
5.564006E+3   1.000307E+2   1.000307E+2   2.000000E+0   2.000000E+0   9.000000E+1   3.000000E+0   3.000000E+0   -6.761313E-2   8.929601E-2   -9.995915E-5   -8.370437E-6   8.370437E-6   -9.995915E-5   1.003090E-4   -1.752133E+2   -8.521330E+1   
5.585594E+3   1.000484E+2   1.000484E+2   5.000000E+0   5.000000E+0   9.000000E+1   5.000000E+0   5.000000E+0   -6.599450E-2   9.020598E-2   -9.955108E-5   -1.016253E-5   1.016253E-5   -9.955108E-5   1.000685E-4   -1.741712E+2   -8.417123E+1   
5.607347E+3   1.000844E+2   1.000844E+2   6.000000E+0   6.000000E+0   9.000000E+1   8.000000E+0   8.000000E+0   -6.687623E-2   8.956232E-2   -9.967700E-5   -9.089573E-6   9.089573E-6   -9.967700E-5   1.000906E-4   -1.747896E+2   -8.478959E+1   
5.628890E+3   1.000494E+2   1.000494E+2   8.000000E+0   8.000000E+0   9.000000E+1   9.000000E+0   9.000000E+0   -6.722597E-2   9.022134E-2   -1.003224E-4   -9.261749E-6   9.261749E-6   -1.003224E-4   1.007491E-4   -1.747254E+2   -8.472542E+1   
5.650767E+3   9.994451E+1   9.994451E+1   1.000000E+1   1.000000E+1   9.000000E+1   1.100000E+1   1.100000E+1   -6.721982E-2   8.850264E-2   -9.919927E-5   -8.142657E-6   8.142657E-6   -9.919927E-5   9.953290E-5   -1.753075E+2   -8.530746E+1   
5.672595E+3   1.000380E+2   1.000380E+2   1.200000E+1   1.200000E+1   9.000000E+1   1.300000E+1   1.300000E+1   -6.702839E-2   9.035877E-2   -1.002898E-4   -9.497733E-6   9.497733E-6   -1.002898E-4   1.007385E-4   -1.745901E+2   -8.459006E+1   
5.694520E+3   1.000662E+2   1.000662E+2   1.500000E+1   1.500000E+1   9.000000E+1   1.500000E+1   1.500000E+1   -6.626632E-2   8.984090E-2   -9.948137E-5   -9.722812E-6   9.722812E-6   -9.948137E-5   9.995537E-5   -1.744179E+2   -8.441793E+1   
5.716548E+3   1.000387E+2   1.000387E+2   1.600000E+1   1.600000E+1   9.000000E+1   1.700000E+1   1.700000E+1   -6.681120E-2   9.000412E-2   -9.992454E-5   -9.426512E-6   9.426512E-6   -9.992454E-5   1.003682E-4   -1.746109E+2   -8.461088E+1   
5.738435E+3   1.000687E+2   1.000687E+2   1.800000E+1   1.800000E+1   9.000000E+1   1.900000E+1   1.900000E+1   -6.717014E-2   9.062751E-2   -1.005525E-4   -9.568582E-6   9.568582E-6   -1.005525E-4   1.010067E-4   -1.745641E+2   -8.456410E+1   
5.760310E+3   1.000530E+2   1.000530E+2   2.000000E+1   2.000000E+1   9.000000E+1   2.100000E+1   2.100000E+1   -6.689280E-2   8.970283E-2   -9.977876E-5   -9.169183E-6   9.169183E-6   -9.977876E-5   1.001992E-4   -1.747495E+2   -8.474954E+1   
5.782188E+3   1.000146E+2   1.000146E+2   2.200000E+1   2.200000E+1   9.000000E+1   2.300000E+1   2.300000E+1   -6.761314E-2   9.042809E-2   -1.006965E-4   -9.110555E-6   9.110555E-6   -1.006965E-4   1.011078E-4   -1.748302E+2   -8.483022E+1   
5.804026E+3   1.000366E+2   1.000366E+2   2.400000E+1   2.400000E+1   9.000000E+1   2.500000E+1   2.500000E+1   -6.752786E-2   9.086191E-2   -1.009263E-4   -9.457248E-6   9.457248E-6   -1.009263E-4   1.013684E-4   -1.746468E+2   -8.464676E+1   
5.825907E+3   1.000217E+2   1.000217E+2   2.600000E+1   2.600000E+1   9.000000E+1   2.700000E+1   2.700000E+1   -6.690138E-2   8.946046E-2   -9.962621E-5   -9.004381E-6   9.004381E-6   -9.962621E-5   1.000323E-4   -1.748355E+2   -8.483555E+1   
5.847834E+3   1.000124E+2   1.000124E+2   2.800000E+1   2.800000E+1   9.000000E+1   2.900000E+1   2.900000E+1   -6.710939E-2   9.118404E-2   -1.008774E-4   -9.977361E-6   9.977361E-6   -1.008774E-4   1.013696E-4   -1.743515E+2   -8.435148E+1   
5.869750E+3   9.999371E+1   9.999371E+1   3.000000E+1   3.000000E+1   9.000000E+1   3.100000E+1   3.100000E+1   -6.776715E-2   9.020662E-2   -1.006474E-4   -8.851848E-6   8.851848E-6   -1.006474E-4   1.010359E-4   -1.749738E+2   -8.497382E+1   
5.891697E+3   1.000382E+2   1.000382E+2   3.200000E+1   3.200000E+1   9.000000E+1   3.300000E+1   3.300000E+1   -6.821261E-2   8.981208E-2   -1.006659E-4   -8.264437E-6   8.264437E-6   -1.006659E-4   1.010046E-4   -1.753067E+2   -8.530667E+1   
5.913596E+3   1.000554E+2   1.000554E+2   3.400000E+1   3.400000E+1   9.000000E+1   3.500000E+1   3.500000E+1   -6.770578E-2   9.055023E-2   -1.008333E-4   -9.121880E-6   9.121880E-6   -1.008333E-4   1.012450E-4   -1.748308E+2   -8.483081E+1   
5.935472E+3   1.000193E+2   1.000193E+2   3.600000E+1   3.600000E+1   9.000000E+1   3.700000E+1   3.700000E+1   -6.738673E-2   9.088956E-2   -1.008570E-4   -9.579708E-6   9.579708E-6   -1.008570E-4   1.013110E-4   -1.745742E+2   -8.457415E+1   
5.957442E+3   1.000087E+2   1.000087E+2   3.800000E+1   3.800000E+1   9.000000E+1   3.900000E+1   3.900000E+1   -6.766774E-2   9.031888E-2   -1.006591E-4   -8.998771E-6   8.998771E-6   -1.006591E-4   1.010605E-4   -1.748914E+2   -8.489142E+1   
5.979312E+3   1.001117E+2   1.001117E+2   4.000000E+1   4.000000E+1   9.000000E+1   4.100000E+1   4.100000E+1   -6.635468E-2   9.073737E-2   -1.001199E-4   -1.024355E-5   1.024355E-5   -1.001199E-4   1.006425E-4   -1.741582E+2   -8.415823E+1   
6.001201E+3   1.000469E+2   1.000469E+2   4.200000E+1   4.200000E+1   9.000000E+1   4.300000E+1   4.300000E+1   -6.707318E-2   9.117055E-2   -1.008462E-4   -9.995325E-6   9.995325E-6   -1.008462E-4   1.013403E-4   -1.743396E+2   -8.433964E+1   
6.023059E+3   1.000044E+2   1.000044E+2   4.400000E+1   4.400000E+1   9.000000E+1   4.500000E+1   4.500000E+1   -6.730266E-2   9.013849E-2   -1.003159E-4   -9.150860E-6   9.150860E-6   -1.003159E-4   1.007324E-4   -1.747879E+2   -8.478788E+1   
6.044931E+3   1.000232E+2   1.000232E+2   4.600000E+1   4.600000E+1   9.000000E+1   4.700000E+1   4.700000E+1   -6.735359E-2   9.126015E-2   -1.010779E-4   -9.846496E-6   9.846496E-6   -1.010779E-4   1.015564E-4   -1.744361E+2   -8.443609E+1   
6.066831E+3   1.000551E+2   1.000551E+2   4.800000E+1   4.800000E+1   9.000000E+1   4.900000E+1   4.900000E+1   -6.690507E-2   9.055570E-2   -1.003418E-4   -9.717690E-6   9.717690E-6   -1.003418E-4   1.008113E-4   -1.744684E+2   -8.446839E+1   
6.100791E+3   1.000190E+2   1.000190E+2   9.800000E+1   9.800000E+1   9.000000E+1   9.900000E+1   9.900000E+1   -6.817704E-2   9.308195E-2   -1.027735E-4   -1.042849E-5   1.042849E-5   -1.027735E-4   1.033013E-4   -1.742060E+2   -8.420599E+1   
6.123351E+3   1.000727E+2   1.000727E+2   1.480000E+2   1.480000E+2   9.000000E+1   1.490000E+2   1.490000E+2   -6.963062E-2   9.386309E-2   -1.041809E-4   -9.864066E-6   9.864066E-6   -1.041809E-4   1.046469E-4   -1.745912E+2   -8.459124E+1   
6.145531E+3   1.000340E+2   1.000340E+2   1.980000E+2   1.980000E+2   9.000000E+1   1.990000E+2   1.990000E+2   -7.084244E-2   9.547507E-2   -1.059800E-4   -1.002164E-5   1.002164E-5   -1.059800E-4   1.064528E-4   -1.745981E+2   -8.459808E+1   
6.167921E+3   1.000295E+2   1.000295E+2   2.480000E+2   2.480000E+2   9.000000E+1   2.490000E+2   2.490000E+2   -7.048655E-2   9.767914E-2   -1.071955E-4   -1.172582E-5   1.172582E-5   -1.071955E-4   1.078349E-4   -1.737574E+2   -8.375739E+1   
6.190858E+3   1.000284E+2   1.000284E+2   2.980000E+2   2.980000E+2   9.000000E+1   2.990000E+2   2.990000E+2   -7.418465E-2   9.806262E-2   -1.097316E-4   -9.241297E-6   9.241297E-6   -1.097316E-4   1.101200E-4   -1.751861E+2   -8.518606E+1   
6.213040E+3   1.000066E+2   1.000066E+2   3.480000E+2   3.480000E+2   9.000000E+1   3.490000E+2   3.490000E+2   -7.390547E-2   1.002329E-1   -1.109725E-4   -1.086668E-5   1.086668E-5   -1.109725E-4   1.115032E-4   -1.744073E+2   -8.440730E+1   
6.235380E+3   1.000288E+2   1.000288E+2   3.980000E+2   3.980000E+2   9.000000E+1   3.990000E+2   3.990000E+2   -7.494059E-2   1.013006E-1   -1.123078E-4   -1.079905E-5   1.079905E-5   -1.123078E-4   1.128258E-4   -1.745076E+2   -8.450756E+1   
6.258255E+3   1.000317E+2   1.000317E+2   4.480000E+2   4.480000E+2   9.000000E+1   4.490000E+2   4.490000E+2   -7.317099E-2   1.025664E-1   -1.120381E-4   -1.293547E-5   1.293547E-5   -1.120381E-4   1.127824E-4   -1.734140E+2   -8.341402E+1   
6.280376E+3   9.997589E+1   9.997589E+1   4.980000E+2   4.980000E+2   9.000000E+1   4.990000E+2   4.990000E+2   -7.570020E-2   1.039445E-1   -1.144994E-4   -1.196576E-5   1.196576E-5   -1.144994E-4   1.151229E-4   -1.740340E+2   -8.403396E+1   
6.302943E+3   9.995010E+1   9.995010E+1   5.480000E+2   5.480000E+2   9.000000E+1   5.490000E+2   5.490000E+2   -7.768760E-2   1.064007E-1   -1.173277E-4   -1.210159E-5   1.210159E-5   -1.173277E-4   1.179502E-4   -1.741111E+2   -8.411114E+1   
6.326278E+3   1.000301E+2   1.000301E+2   5.980000E+2   5.980000E+2   9.000000E+1   5.980000E+2   5.980000E+2   -7.829689E-2   1.077874E-1   -1.186076E-4   -1.255753E-5   1.255753E-5   -1.186076E-4   1.192705E-4   -1.739563E+2   -8.395635E+1   
6.348903E+3   9.996160E+1   9.996160E+1   6.470000E+2   6.470000E+2   9.000000E+1   6.480000E+2   6.480000E+2   -7.931298E-2   1.081396E-1   -1.194651E-4   -1.203625E-5   1.203625E-5   -1.194651E-4   1.200699E-4   -1.742468E+2   -8.424680E+1   
6.371778E+3   1.000241E+2   1.000241E+2   6.970000E+2   6.970000E+2   9.000000E+1   6.980000E+2   6.980000E+2   -8.066102E-2   1.107240E-1   -1.219818E-4   -1.272882E-5   1.272882E-5   -1.219818E-4   1.226441E-4   -1.740427E+2   -8.404273E+1   
6.395080E+3   1.000239E+2   1.000239E+2   7.470000E+2   7.470000E+2   9.000000E+1   7.480000E+2   7.480000E+2   -8.102735E-2   1.117996E-1   -1.229088E-4   -1.316108E-5   1.316108E-5   -1.229088E-4   1.236114E-4   -1.738881E+2   -8.388805E+1   
6.417696E+3   1.000686E+2   1.000686E+2   7.970000E+2   7.970000E+2   9.000000E+1   7.980000E+2   7.980000E+2   -8.250238E-2   1.129378E-1   -1.245620E-4   -1.281422E-5   1.281422E-5   -1.245620E-4   1.252194E-4   -1.741264E+2   -8.412640E+1   
6.440338E+3   1.000181E+2   1.000181E+2   8.470000E+2   8.470000E+2   9.000000E+1   8.480000E+2   8.480000E+2   -8.325833E-2   1.144540E-1   -1.260169E-4   -1.324634E-5   1.324634E-5   -1.260169E-4   1.267111E-4   -1.739994E+2   -8.399936E+1   
6.463620E+3   1.000085E+2   1.000085E+2   8.980000E+2   8.980000E+2   9.000000E+1   8.980000E+2   8.980000E+2   -8.362343E-2   1.155560E-1   -1.269603E-4   -1.369674E-5   1.369674E-5   -1.269603E-4   1.276970E-4   -1.738426E+2   -8.384262E+1   
6.486210E+3   1.000636E+2   1.000636E+2   9.470000E+2   9.470000E+2   9.000000E+1   9.480000E+2   9.480000E+2   -8.625509E-2   1.180514E-1   -1.302126E-4   -1.338174E-5   1.338174E-5   -1.302126E-4   1.308984E-4   -1.741324E+2   -8.413240E+1   
6.508761E+3   9.997650E+1   9.997650E+1   9.970000E+2   9.970000E+2   9.000000E+1   9.980000E+2   9.980000E+2   -8.576299E-2   1.206586E-1   -1.316063E-4   -1.545019E-5   1.545019E-5   -1.316063E-4   1.325101E-4   -1.733043E+2   -8.330430E+1   
6.532306E+3   9.998531E+1   9.998531E+1   1.047000E+3   1.047000E+3   9.000000E+1   1.048000E+3   1.048000E+3   -8.681835E-2   1.206794E-1   -1.322724E-4   -1.468325E-5   1.468325E-5   -1.322724E-4   1.330849E-4   -1.736657E+2   -8.366566E+1   
6.555091E+3   1.000319E+2   1.000319E+2   1.098000E+3   1.098000E+3   9.000000E+1   1.098000E+3   1.098000E+3   -8.715644E-2   1.228834E-1   -1.339168E-4   -1.587408E-5   1.587408E-5   -1.339168E-4   1.348544E-4   -1.732399E+2   -8.323988E+1   
6.577926E+3   9.997311E+1   9.997311E+1   1.148000E+3   1.148000E+3   9.000000E+1   1.148000E+3   1.148000E+3   -8.936415E-2   1.238590E-1   -1.359172E-4   -1.487902E-5   1.487902E-5   -1.359172E-4   1.367291E-4   -1.737526E+2   -8.375264E+1   
6.601194E+3   1.000155E+2   1.000155E+2   1.198000E+3   1.198000E+3   9.000000E+1   1.199000E+3   1.199000E+3   -9.008695E-2   1.260207E-1   -1.377719E-4   -1.575766E-5   1.575766E-5   -1.377719E-4   1.386701E-4   -1.734752E+2   -8.347515E+1   
6.624035E+3   1.000664E+2   1.000664E+2   1.248000E+3   1.248000E+3   9.000000E+1   1.248000E+3   1.248000E+3   -9.160440E-2   1.265214E-1   -1.390361E-4   -1.496262E-5   1.496262E-5   -1.390361E-4   1.398389E-4   -1.738577E+2   -8.385765E+1   
6.646610E+3   1.000505E+2   1.000505E+2   1.298000E+3   1.298000E+3   9.000000E+1   1.298000E+3   1.298000E+3   -9.180991E-2   1.282014E-1   -1.402574E-4   -1.590897E-5   1.590897E-5   -1.402574E-4   1.411567E-4   -1.735288E+2   -8.352877E+1   
6.670110E+3   1.000344E+2   1.000344E+2   1.348000E+3   1.348000E+3   9.000000E+1   1.349000E+3   1.349000E+3   -9.263218E-2   1.295132E-1   -1.416201E-4   -1.615843E-5   1.615843E-5   -1.416201E-4   1.425390E-4   -1.734909E+2   -8.349087E+1   
6.692661E+3   1.000224E+2   1.000224E+2   1.398000E+3   1.398000E+3   9.000000E+1   1.399000E+3   1.399000E+3   -9.379253E-2   1.308398E-1   -1.432015E-4   -1.616748E-5   1.616748E-5   -1.432015E-4   1.441112E-4   -1.735586E+2   -8.355857E+1   
6.715642E+3   1.000033E+2   1.000033E+2   1.448000E+3   1.448000E+3   9.000000E+1   1.449000E+3   1.449000E+3   -9.431044E-2   1.334248E-1   -1.452053E-4   -1.747444E-5   1.747444E-5   -1.452053E-4   1.462530E-4   -1.731379E+2   -8.313785E+1   
6.738734E+3   1.000410E+2   1.000410E+2   1.498000E+3   1.498000E+3   9.000000E+1   1.499000E+3   1.499000E+3   -9.540939E-2   1.343458E-1   -1.464845E-4   -1.726373E-5   1.726373E-5   -1.464845E-4   1.474983E-4   -1.732785E+2   -8.327849E+1   
6.761345E+3   1.000392E+2   1.000392E+2   1.548000E+3   1.548000E+3   9.000000E+1   1.549000E+3   1.549000E+3   -9.551067E-2   1.365449E-1   -1.479794E-4   -1.862652E-5   1.862652E-5   -1.479794E-4   1.491471E-4   -1.728258E+2   -8.282577E+1   
6.783905E+3   1.000221E+2   1.000221E+2   1.598000E+3   1.598000E+3   9.000000E+1   1.599000E+3   1.599000E+3   -9.904501E-2   1.374567E-1   -1.507583E-4   -1.660852E-5   1.660852E-5   -1.507583E-4   1.516704E-4   -1.737133E+2   -8.371327E+1   
6.806983E+3   1.000230E+2   1.000230E+2   1.648000E+3   1.648000E+3   9.000000E+1   1.649000E+3   1.649000E+3   -9.981936E-2   1.381930E-1   -1.517166E-4   -1.651717E-5   1.651717E-5   -1.517166E-4   1.526131E-4   -1.737868E+2   -8.378676E+1   
6.829564E+3   1.000466E+2   1.000466E+2   1.698000E+3   1.698000E+3   9.000000E+1   1.699000E+3   1.699000E+3   -9.871917E-2   1.396410E-1   -1.519795E-4   -1.827759E-5   1.827759E-5   -1.519795E-4   1.530747E-4   -1.731423E+2   -8.314234E+1   
6.852141E+3   1.000619E+2   1.000619E+2   1.748000E+3   1.748000E+3   9.000000E+1   1.749000E+3   1.749000E+3   -1.001372E-1   1.415020E-1   -1.540683E-4   -1.844546E-5   1.844546E-5   -1.540683E-4   1.551685E-4   -1.731729E+2   -8.317289E+1   
6.874921E+3   9.999441E+1   9.999441E+1   1.798000E+3   1.798000E+3   9.000000E+1   1.799000E+3   1.799000E+3   -1.009048E-1   1.435483E-1   -1.558756E-4   -1.921553E-5   1.921553E-5   -1.558756E-4   1.570555E-4   -1.729723E+2   -8.297233E+1   
6.897495E+3   1.000634E+2   1.000634E+2   1.848000E+3   1.848000E+3   9.000000E+1   1.849000E+3   1.849000E+3   -1.020724E-1   1.446129E-1   -1.572908E-4   -1.904789E-5   1.904789E-5   -1.572908E-4   1.584400E-4   -1.730951E+2   -8.309511E+1   
6.920073E+3   1.000081E+2   1.000081E+2   1.898000E+3   1.898000E+3   9.000000E+1   1.899000E+3   1.899000E+3   -1.031757E-1   1.466635E-1   -1.593084E-4   -1.957254E-5   1.957254E-5   -1.593084E-4   1.605063E-4   -1.729958E+2   -8.299578E+1   
6.942846E+3   1.000342E+2   1.000342E+2   1.948000E+3   1.948000E+3   9.000000E+1   1.949000E+3   1.949000E+3   -1.036653E-1   1.474710E-1   -1.601370E-4   -1.973828E-5   1.973828E-5   -1.601370E-4   1.613489E-4   -1.729732E+2   -8.297324E+1   
6.965392E+3   1.000460E+2   1.000460E+2   1.998000E+3   1.998000E+3   9.000000E+1   1.999000E+3   1.999000E+3   -1.046225E-1   1.490411E-1   -1.617514E-4   -2.005684E-5   2.005684E-5   -1.617514E-4   1.629902E-4   -1.729315E+2   -8.293152E+1   
7.003334E+3   1.000427E+2   1.000427E+2   2.498000E+3   2.498000E+3   9.000000E+1   2.499000E+3   2.499000E+3   -1.165739E-1   1.655853E-1   -1.799154E-4   -2.203327E-5   2.203327E-5   -1.799154E-4   1.812595E-4   -1.730181E+2   -8.301806E+1   
7.029780E+3   9.998919E+1   9.998919E+1   2.998000E+3   2.998000E+3   9.000000E+1   2.999000E+3   2.999000E+3   -1.265852E-1   1.811133E-1   -1.962180E-4   -2.478042E-5   2.478042E-5   -1.962180E-4   1.977766E-4   -1.728022E+2   -8.280221E+1   
7.055724E+3   1.000566E+2   1.000566E+2   3.498000E+3   3.498000E+3   9.000000E+1   3.499000E+3   3.499000E+3   -1.364289E-1   1.974715E-1   -2.129579E-4   -2.819424E-5   2.819424E-5   -2.129579E-4   2.148161E-4   -1.724583E+2   -8.245827E+1   
7.081587E+3   1.000160E+2   1.000160E+2   3.998000E+3   3.998000E+3   9.000000E+1   3.999000E+3   3.999000E+3   -1.477594E-1   2.136512E-1   -2.305005E-4   -3.039167E-5   3.039167E-5   -2.305005E-4   2.324955E-4   -1.724888E+2   -8.248883E+1   
7.108229E+3   9.997360E+1   9.997360E+1   4.498000E+3   4.498000E+3   9.000000E+1   4.498000E+3   4.498000E+3   -1.544002E-1   2.248411E-1   -2.418941E-4   -3.279557E-5   3.279557E-5   -2.418941E-4   2.441071E-4   -1.722790E+2   -8.227902E+1   
7.134379E+3   9.998959E+1   9.998959E+1   4.997000E+3   4.997000E+3   9.000000E+1   4.998000E+3   4.998000E+3   -1.549708E-1   2.277556E-1   -2.441451E-4   -3.427896E-5   3.427896E-5   -2.441451E-4   2.465398E-4   -1.720077E+2   -8.200768E+1   
7.160072E+3   1.000061E+2   1.000061E+2   5.498000E+3   5.498000E+3   9.000000E+1   5.499000E+3   5.499000E+3   -1.472673E-1   2.222309E-1   -2.357842E-4   -3.636484E-5   3.636484E-5   -2.357842E-4   2.385719E-4   -1.712324E+2   -8.123239E+1   
7.186516E+3   1.000218E+2   1.000218E+2   5.998000E+3   5.998000E+3   9.000000E+1   5.999000E+3   5.999000E+3   -1.301673E-1   2.030374E-1   -2.127116E-4   -3.646434E-5   3.646434E-5   -2.127116E-4   2.158144E-4   -1.702726E+2   -8.027255E+1   
7.212660E+3   9.995870E+1   9.995870E+1   6.498000E+3   6.498000E+3   9.000000E+1   6.498000E+3   6.498000E+3   -1.207046E-1   1.915245E-1   -1.993631E-4   -3.593648E-5   3.593648E-5   -1.993631E-4   2.025761E-4   -1.697818E+2   -7.978180E+1   
7.238815E+3   9.999371E+1   9.999371E+1   6.997000E+3   6.997000E+3   9.000000E+1   6.998000E+3   6.998000E+3   -1.084562E-1   1.815189E-1   -1.852740E-4   -3.845435E-5   3.845435E-5   -1.852740E-4   1.892226E-4   -1.682745E+2   -7.827452E+1   
7.264545E+3   1.000365E+2   1.000365E+2   7.498000E+3   7.498000E+3   9.000000E+1   7.499000E+3   7.499000E+3   -1.085065E-1   1.818741E-1   -1.855365E-4   -3.864938E-5   3.864938E-5   -1.855365E-4   1.895193E-4   -1.682329E+2   -7.823291E+1   
7.290480E+3   1.000227E+2   1.000227E+2   7.999000E+3   7.999000E+3   9.000000E+1   8.000000E+3   8.000000E+3   -1.121021E-1   1.863007E-1   -1.906424E-4   -3.888391E-5   3.888391E-5   -1.906424E-4   1.945674E-4   -1.684719E+2   -7.847193E+1   
7.316859E+3   9.999981E+1   9.999981E+1   8.498000E+3   8.498000E+3   9.000000E+1   8.498000E+3   8.498000E+3   -1.201572E-1   2.006714E-1   -2.049820E-4   -4.232126E-5   4.232126E-5   -2.049820E-4   2.093053E-4   -1.683344E+2   -7.833444E+1   
7.343311E+3   1.000042E+2   1.000042E+2   8.998000E+3   8.998000E+3   9.000000E+1   8.999000E+3   8.999000E+3   -1.351251E-1   2.195668E-1   -2.265421E-4   -4.360385E-5   4.360385E-5   -2.265421E-4   2.307003E-4   -1.691052E+2   -7.910519E+1   
7.369413E+3   9.998760E+1   9.998760E+1   9.498000E+3   9.498000E+3   9.000000E+1   9.499000E+3   9.499000E+3   -1.448093E-1   2.343946E-1   -2.421866E-4   -4.613515E-5   4.613515E-5   -2.421866E-4   2.465417E-4   -1.692147E+2   -7.921471E+1   
7.394860E+3   1.000236E+2   1.000236E+2   9.998000E+3   9.998000E+3   9.000000E+1   9.999000E+3   9.999000E+3   -1.598108E-1   2.553941E-1   -2.651380E-4   -4.876841E-5   4.876841E-5   -2.651380E-4   2.695858E-4   -1.695777E+2   -7.957774E+1   
@@END Data.
@Time at end of measurement: 17:18:06
@NO Instrument  Changes.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   -9499.000      -9998.000      249.500        Coercive Field: Field at which M//H changes sign
Ms  emu                                 3.207E-4       -3.584E-4      3.395E-4       Saturation Magnetization: maximum M measured
Mr emu                                  -9.942E-5      1.332E-4       1.163E-4       Remanent Magnetization: M at H=0        
S                                       0.310          0.372          0.341          Squareness: Mr/Ms                       
S*                                      1.273          1.223          1.248          1-(Mr/Hc)(1/slope at Hc)                
                                                                                                                             

@END Measurement parameters
